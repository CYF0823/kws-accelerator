module Memory(
  input         clock,
  input  [11:0] io_rdAddr,
  output [15:0] io_rdData,
  input         io_wrEna,
  input  [15:0] io_wrData,
  input  [11:0] io_wrAddr
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] mem [0:3199]; // @[Memory.scala 13:24]
  wire [15:0] mem_io_rdData_MPORT_data; // @[Memory.scala 13:24]
  wire [11:0] mem_io_rdData_MPORT_addr; // @[Memory.scala 13:24]
  wire [15:0] mem_MPORT_data; // @[Memory.scala 13:24]
  wire [11:0] mem_MPORT_addr; // @[Memory.scala 13:24]
  wire  mem_MPORT_mask; // @[Memory.scala 13:24]
  wire  mem_MPORT_en; // @[Memory.scala 13:24]
  reg [11:0] mem_io_rdData_MPORT_addr_pipe_0;
  assign mem_io_rdData_MPORT_addr = mem_io_rdData_MPORT_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_io_rdData_MPORT_data = mem[mem_io_rdData_MPORT_addr]; // @[Memory.scala 13:24]
  `else
  assign mem_io_rdData_MPORT_data = mem_io_rdData_MPORT_addr >= 12'hc80 ? _RAND_1[15:0] : mem[mem_io_rdData_MPORT_addr]; // @[Memory.scala 13:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem_MPORT_data = io_wrData;
  assign mem_MPORT_addr = io_wrAddr;
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = io_wrEna;
  assign io_rdData = mem_io_rdData_MPORT_data; // @[Memory.scala 15:13]
  always @(posedge clock) begin
    if(mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data; // @[Memory.scala 13:24]
    end
    mem_io_rdData_MPORT_addr_pipe_0 <= io_rdAddr;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3200; initvar = initvar+1)
    mem[initvar] = _RAND_0[15:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  mem_io_rdData_MPORT_addr_pipe_0 = _RAND_2[11:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MulAddRecFNToRaw_preMul(
  input  [16:0] io_a,
  input  [16:0] io_b,
  input  [16:0] io_c,
  output [10:0] io_mulAddA,
  output [10:0] io_mulAddB,
  output [21:0] io_mulAddC,
  output        io_toPostMul_isSigNaNAny,
  output        io_toPostMul_isNaNAOrB,
  output        io_toPostMul_isInfA,
  output        io_toPostMul_isZeroA,
  output        io_toPostMul_isInfB,
  output        io_toPostMul_isZeroB,
  output        io_toPostMul_signProd,
  output        io_toPostMul_isNaNC,
  output        io_toPostMul_isInfC,
  output        io_toPostMul_isZeroC,
  output [6:0]  io_toPostMul_sExpSum,
  output        io_toPostMul_doSubMags,
  output        io_toPostMul_CIsDominant,
  output [3:0]  io_toPostMul_CDom_CAlignDist,
  output [12:0] io_toPostMul_highAlignedSigC,
  output        io_toPostMul_bit0AlignedSigC
);
  wire [5:0] rawA_exp = io_a[15:10]; // @[rawFloatFromRecFN.scala 50:21]
  wire  rawA_isZero = rawA_exp[5:3] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  wire  rawA_isSpecial = rawA_exp[5:4] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawA__isNaN = rawA_isSpecial & rawA_exp[3]; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawA__sign = io_a[16]; // @[rawFloatFromRecFN.scala 58:25]
  wire [6:0] rawA__sExp = {1'b0,$signed(rawA_exp)}; // @[rawFloatFromRecFN.scala 59:27]
  wire  rawA_out_sig_hi_lo = ~rawA_isZero; // @[rawFloatFromRecFN.scala 60:39]
  wire [9:0] rawA_out_sig_lo = io_a[9:0]; // @[rawFloatFromRecFN.scala 60:51]
  wire [11:0] rawA__sig = {1'h0,rawA_out_sig_hi_lo,rawA_out_sig_lo}; // @[Cat.scala 30:58]
  wire [5:0] rawB_exp = io_b[15:10]; // @[rawFloatFromRecFN.scala 50:21]
  wire  rawB_isZero = rawB_exp[5:3] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  wire  rawB_isSpecial = rawB_exp[5:4] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawB__isNaN = rawB_isSpecial & rawB_exp[3]; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawB__sign = io_b[16]; // @[rawFloatFromRecFN.scala 58:25]
  wire [6:0] rawB__sExp = {1'b0,$signed(rawB_exp)}; // @[rawFloatFromRecFN.scala 59:27]
  wire  rawB_out_sig_hi_lo = ~rawB_isZero; // @[rawFloatFromRecFN.scala 60:39]
  wire [9:0] rawB_out_sig_lo = io_b[9:0]; // @[rawFloatFromRecFN.scala 60:51]
  wire [11:0] rawB__sig = {1'h0,rawB_out_sig_hi_lo,rawB_out_sig_lo}; // @[Cat.scala 30:58]
  wire [5:0] rawC_exp = io_c[15:10]; // @[rawFloatFromRecFN.scala 50:21]
  wire  rawC_isZero = rawC_exp[5:3] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  wire  rawC_isSpecial = rawC_exp[5:4] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawC__isNaN = rawC_isSpecial & rawC_exp[3]; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawC__sign = io_c[16]; // @[rawFloatFromRecFN.scala 58:25]
  wire [6:0] rawC__sExp = {1'b0,$signed(rawC_exp)}; // @[rawFloatFromRecFN.scala 59:27]
  wire  rawC_out_sig_hi_lo = ~rawC_isZero; // @[rawFloatFromRecFN.scala 60:39]
  wire [9:0] rawC_out_sig_lo = io_c[9:0]; // @[rawFloatFromRecFN.scala 60:51]
  wire [11:0] rawC__sig = {1'h0,rawC_out_sig_hi_lo,rawC_out_sig_lo}; // @[Cat.scala 30:58]
  wire  signProd = rawA__sign ^ rawB__sign; // @[MulAddRecFN.scala 100:30]
  wire [7:0] _sExpAlignedProd_T = $signed(rawA__sExp) + $signed(rawB__sExp); // @[MulAddRecFN.scala 103:19]
  wire [7:0] sExpAlignedProd = $signed(_sExpAlignedProd_T) - 8'sh12; // @[MulAddRecFN.scala 103:32]
  wire  doSubMags = signProd ^ rawC__sign; // @[MulAddRecFN.scala 105:30]
  wire [7:0] _GEN_0 = {{1{rawC__sExp[6]}},rawC__sExp}; // @[MulAddRecFN.scala 109:42]
  wire [7:0] sNatCAlignDist = $signed(sExpAlignedProd) - $signed(_GEN_0); // @[MulAddRecFN.scala 109:42]
  wire [6:0] posNatCAlignDist = sNatCAlignDist[6:0]; // @[MulAddRecFN.scala 110:42]
  wire  isMinCAlign = rawA_isZero | rawB_isZero | $signed(sNatCAlignDist) < 8'sh0; // @[MulAddRecFN.scala 111:50]
  wire  CIsDominant = rawC_out_sig_hi_lo & (isMinCAlign | posNatCAlignDist <= 7'hb); // @[MulAddRecFN.scala 113:23]
  wire [5:0] _CAlignDist_T_2 = posNatCAlignDist < 7'h23 ? posNatCAlignDist[5:0] : 6'h23; // @[MulAddRecFN.scala 117:16]
  wire [5:0] CAlignDist = isMinCAlign ? 6'h0 : _CAlignDist_T_2; // @[MulAddRecFN.scala 115:12]
  wire [11:0] _mainAlignedSigC_T = ~rawC__sig; // @[MulAddRecFN.scala 123:28]
  wire [11:0] mainAlignedSigC_hi = doSubMags ? _mainAlignedSigC_T : rawC__sig; // @[MulAddRecFN.scala 123:16]
  wire [26:0] mainAlignedSigC_lo = doSubMags ? 27'h7ffffff : 27'h0; // @[Bitwise.scala 72:12]
  wire [38:0] _mainAlignedSigC_T_3 = {mainAlignedSigC_hi,mainAlignedSigC_lo}; // @[MulAddRecFN.scala 125:11]
  wire [38:0] mainAlignedSigC = $signed(_mainAlignedSigC_T_3) >>> CAlignDist; // @[MulAddRecFN.scala 125:17]
  wire  reduced4CExtra_reducedVec_0 = |rawC__sig[3:0]; // @[primitives.scala 121:54]
  wire  reduced4CExtra_reducedVec_1 = |rawC__sig[7:4]; // @[primitives.scala 121:54]
  wire  reduced4CExtra_reducedVec_2 = |rawC__sig[11:8]; // @[primitives.scala 124:57]
  wire [2:0] _reduced4CExtra_T_1 = {reduced4CExtra_reducedVec_2,reduced4CExtra_reducedVec_1,reduced4CExtra_reducedVec_0}
    ; // @[primitives.scala 125:20]
  wire [16:0] reduced4CExtra_shift = 17'sh10000 >>> CAlignDist[5:2]; // @[primitives.scala 77:58]
  wire  reduced4CExtra_hi_1 = reduced4CExtra_shift[8]; // @[Bitwise.scala 109:18]
  wire  reduced4CExtra_lo = reduced4CExtra_shift[9]; // @[Bitwise.scala 109:44]
  wire [1:0] _reduced4CExtra_T_4 = {reduced4CExtra_hi_1,reduced4CExtra_lo}; // @[Cat.scala 30:58]
  wire [2:0] _GEN_1 = {{1'd0}, _reduced4CExtra_T_4}; // @[MulAddRecFN.scala 127:68]
  wire [2:0] _reduced4CExtra_T_5 = _reduced4CExtra_T_1 & _GEN_1; // @[MulAddRecFN.scala 127:68]
  wire  reduced4CExtra = |_reduced4CExtra_T_5; // @[MulAddRecFN.scala 135:11]
  wire  _alignedSigC_T_4 = &mainAlignedSigC[2:0] & ~reduced4CExtra; // @[MulAddRecFN.scala 139:44]
  wire  _alignedSigC_T_7 = |mainAlignedSigC[2:0] | reduced4CExtra; // @[MulAddRecFN.scala 140:44]
  wire  alignedSigC_lo = doSubMags ? _alignedSigC_T_4 : _alignedSigC_T_7; // @[MulAddRecFN.scala 138:16]
  wire [35:0] alignedSigC_hi = mainAlignedSigC[38:3]; // @[Cat.scala 30:58]
  wire [36:0] alignedSigC = {alignedSigC_hi,alignedSigC_lo}; // @[Cat.scala 30:58]
  wire  _io_toPostMul_isSigNaNAny_T_2 = rawA__isNaN & ~rawA__sig[9]; // @[common.scala 81:46]
  wire  _io_toPostMul_isSigNaNAny_T_5 = rawB__isNaN & ~rawB__sig[9]; // @[common.scala 81:46]
  wire  _io_toPostMul_isSigNaNAny_T_9 = rawC__isNaN & ~rawC__sig[9]; // @[common.scala 81:46]
  wire [7:0] _io_toPostMul_sExpSum_T_2 = $signed(sExpAlignedProd) - 8'shb; // @[MulAddRecFN.scala 163:53]
  wire [7:0] _io_toPostMul_sExpSum_T_3 = CIsDominant ? $signed({{1{rawC__sExp[6]}},rawC__sExp}) : $signed(
    _io_toPostMul_sExpSum_T_2); // @[MulAddRecFN.scala 163:12]
  assign io_mulAddA = rawA__sig[10:0]; // @[MulAddRecFN.scala 146:16]
  assign io_mulAddB = rawB__sig[10:0]; // @[MulAddRecFN.scala 147:16]
  assign io_mulAddC = alignedSigC[22:1]; // @[MulAddRecFN.scala 148:30]
  assign io_toPostMul_isSigNaNAny = _io_toPostMul_isSigNaNAny_T_2 | _io_toPostMul_isSigNaNAny_T_5 |
    _io_toPostMul_isSigNaNAny_T_9; // @[MulAddRecFN.scala 151:58]
  assign io_toPostMul_isNaNAOrB = rawA__isNaN | rawB__isNaN; // @[MulAddRecFN.scala 153:42]
  assign io_toPostMul_isInfA = rawA_isSpecial & ~rawA_exp[3]; // @[rawFloatFromRecFN.scala 56:33]
  assign io_toPostMul_isZeroA = rawA_exp[5:3] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign io_toPostMul_isInfB = rawB_isSpecial & ~rawB_exp[3]; // @[rawFloatFromRecFN.scala 56:33]
  assign io_toPostMul_isZeroB = rawB_exp[5:3] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign io_toPostMul_signProd = rawA__sign ^ rawB__sign; // @[MulAddRecFN.scala 100:30]
  assign io_toPostMul_isNaNC = rawC_isSpecial & rawC_exp[3]; // @[rawFloatFromRecFN.scala 55:33]
  assign io_toPostMul_isInfC = rawC_isSpecial & ~rawC_exp[3]; // @[rawFloatFromRecFN.scala 56:33]
  assign io_toPostMul_isZeroC = rawC_exp[5:3] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  assign io_toPostMul_sExpSum = _io_toPostMul_sExpSum_T_3[6:0]; // @[MulAddRecFN.scala 162:28]
  assign io_toPostMul_doSubMags = signProd ^ rawC__sign; // @[MulAddRecFN.scala 105:30]
  assign io_toPostMul_CIsDominant = rawC_out_sig_hi_lo & (isMinCAlign | posNatCAlignDist <= 7'hb); // @[MulAddRecFN.scala 113:23]
  assign io_toPostMul_CDom_CAlignDist = CAlignDist[3:0]; // @[MulAddRecFN.scala 166:47]
  assign io_toPostMul_highAlignedSigC = alignedSigC[35:23]; // @[MulAddRecFN.scala 168:20]
  assign io_toPostMul_bit0AlignedSigC = alignedSigC[0]; // @[MulAddRecFN.scala 169:48]
endmodule
module MulAddRecFNToRaw_postMul(
  input         io_fromPreMul_isSigNaNAny,
  input         io_fromPreMul_isNaNAOrB,
  input         io_fromPreMul_isInfA,
  input         io_fromPreMul_isZeroA,
  input         io_fromPreMul_isInfB,
  input         io_fromPreMul_isZeroB,
  input         io_fromPreMul_signProd,
  input         io_fromPreMul_isNaNC,
  input         io_fromPreMul_isInfC,
  input         io_fromPreMul_isZeroC,
  input  [6:0]  io_fromPreMul_sExpSum,
  input         io_fromPreMul_doSubMags,
  input         io_fromPreMul_CIsDominant,
  input  [3:0]  io_fromPreMul_CDom_CAlignDist,
  input  [12:0] io_fromPreMul_highAlignedSigC,
  input         io_fromPreMul_bit0AlignedSigC,
  input  [22:0] io_mulAddResult,
  output        io_invalidExc,
  output        io_rawOut_isNaN,
  output        io_rawOut_isInf,
  output        io_rawOut_isZero,
  output        io_rawOut_sign,
  output [6:0]  io_rawOut_sExp,
  output [13:0] io_rawOut_sig
);
  wire  CDom_sign = io_fromPreMul_signProd ^ io_fromPreMul_doSubMags; // @[MulAddRecFN.scala 194:42]
  wire [12:0] _sigSum_T_2 = io_fromPreMul_highAlignedSigC + 13'h1; // @[MulAddRecFN.scala 197:47]
  wire [12:0] sigSum_hi_hi = io_mulAddResult[22] ? _sigSum_T_2 : io_fromPreMul_highAlignedSigC; // @[MulAddRecFN.scala 196:16]
  wire [21:0] sigSum_hi_lo = io_mulAddResult[21:0]; // @[MulAddRecFN.scala 200:28]
  wire [35:0] sigSum = {sigSum_hi_hi,sigSum_hi_lo,io_fromPreMul_bit0AlignedSigC}; // @[Cat.scala 30:58]
  wire [1:0] _CDom_sExp_T = {1'b0,$signed(io_fromPreMul_doSubMags)}; // @[MulAddRecFN.scala 207:69]
  wire [6:0] _GEN_0 = {{5{_CDom_sExp_T[1]}},_CDom_sExp_T}; // @[MulAddRecFN.scala 207:43]
  wire [6:0] CDom_sExp = $signed(io_fromPreMul_sExpSum) - $signed(_GEN_0); // @[MulAddRecFN.scala 207:43]
  wire [23:0] _CDom_absSigSum_T_1 = ~sigSum[35:12]; // @[MulAddRecFN.scala 210:13]
  wire [1:0] CDom_absSigSum_hi_lo = io_fromPreMul_highAlignedSigC[12:11]; // @[MulAddRecFN.scala 213:46]
  wire [20:0] CDom_absSigSum_lo = sigSum[33:13]; // @[MulAddRecFN.scala 214:23]
  wire [23:0] _CDom_absSigSum_T_2 = {1'h0,CDom_absSigSum_hi_lo,CDom_absSigSum_lo}; // @[Cat.scala 30:58]
  wire [23:0] CDom_absSigSum = io_fromPreMul_doSubMags ? _CDom_absSigSum_T_1 : _CDom_absSigSum_T_2; // @[MulAddRecFN.scala 209:12]
  wire [10:0] _CDom_absSigSumExtra_T_1 = ~sigSum[11:1]; // @[MulAddRecFN.scala 219:14]
  wire  _CDom_absSigSumExtra_T_2 = |_CDom_absSigSumExtra_T_1; // @[MulAddRecFN.scala 219:36]
  wire  _CDom_absSigSumExtra_T_4 = |sigSum[12:1]; // @[MulAddRecFN.scala 220:37]
  wire  CDom_absSigSumExtra = io_fromPreMul_doSubMags ? _CDom_absSigSumExtra_T_2 : _CDom_absSigSumExtra_T_4; // @[MulAddRecFN.scala 218:12]
  wire [38:0] _GEN_1 = {{15'd0}, CDom_absSigSum}; // @[MulAddRecFN.scala 223:24]
  wire [38:0] _CDom_mainSig_T = _GEN_1 << io_fromPreMul_CDom_CAlignDist; // @[MulAddRecFN.scala 223:24]
  wire [15:0] CDom_mainSig = _CDom_mainSig_T[23:8]; // @[MulAddRecFN.scala 223:56]
  wire  CDom_reduced4SigExtra_reducedVec_0 = |CDom_absSigSum[3:0]; // @[primitives.scala 121:54]
  wire  CDom_reduced4SigExtra_reducedVec_1 = |CDom_absSigSum[7:4]; // @[primitives.scala 121:54]
  wire  CDom_reduced4SigExtra_reducedVec_2 = |CDom_absSigSum[10:8]; // @[primitives.scala 124:57]
  wire [2:0] _CDom_reduced4SigExtra_T_2 = {CDom_reduced4SigExtra_reducedVec_2,CDom_reduced4SigExtra_reducedVec_1,
    CDom_reduced4SigExtra_reducedVec_0}; // @[primitives.scala 125:20]
  wire [1:0] _CDom_reduced4SigExtra_T_4 = ~io_fromPreMul_CDom_CAlignDist[3:2]; // @[primitives.scala 51:21]
  wire [4:0] CDom_reduced4SigExtra_shift = 5'sh10 >>> _CDom_reduced4SigExtra_T_4; // @[primitives.scala 77:58]
  wire  CDom_reduced4SigExtra_hi_1 = CDom_reduced4SigExtra_shift[1]; // @[Bitwise.scala 109:18]
  wire  CDom_reduced4SigExtra_lo = CDom_reduced4SigExtra_shift[2]; // @[Bitwise.scala 109:44]
  wire [1:0] _CDom_reduced4SigExtra_T_6 = {CDom_reduced4SigExtra_hi_1,CDom_reduced4SigExtra_lo}; // @[Cat.scala 30:58]
  wire [2:0] _GEN_2 = {{1'd0}, _CDom_reduced4SigExtra_T_6}; // @[MulAddRecFN.scala 226:72]
  wire [2:0] _CDom_reduced4SigExtra_T_7 = _CDom_reduced4SigExtra_T_2 & _GEN_2; // @[MulAddRecFN.scala 226:72]
  wire  CDom_reduced4SigExtra = |_CDom_reduced4SigExtra_T_7; // @[MulAddRecFN.scala 227:73]
  wire [12:0] CDom_sig_hi = CDom_mainSig[15:3]; // @[MulAddRecFN.scala 229:25]
  wire  CDom_sig_lo = |CDom_mainSig[2:0] | CDom_reduced4SigExtra | CDom_absSigSumExtra; // @[MulAddRecFN.scala 230:61]
  wire [13:0] CDom_sig = {CDom_sig_hi,CDom_sig_lo}; // @[Cat.scala 30:58]
  wire  notCDom_signSigSum = sigSum[25]; // @[MulAddRecFN.scala 236:36]
  wire [24:0] _notCDom_absSigSum_T_1 = ~sigSum[24:0]; // @[MulAddRecFN.scala 239:13]
  wire [24:0] _GEN_3 = {{24'd0}, io_fromPreMul_doSubMags}; // @[MulAddRecFN.scala 240:41]
  wire [24:0] _notCDom_absSigSum_T_4 = sigSum[24:0] + _GEN_3; // @[MulAddRecFN.scala 240:41]
  wire [24:0] notCDom_absSigSum = notCDom_signSigSum ? _notCDom_absSigSum_T_1 : _notCDom_absSigSum_T_4; // @[MulAddRecFN.scala 238:12]
  wire  notCDom_reduced2AbsSigSum_reducedVec_0 = |notCDom_absSigSum[1:0]; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_1 = |notCDom_absSigSum[3:2]; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_2 = |notCDom_absSigSum[5:4]; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_3 = |notCDom_absSigSum[7:6]; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_4 = |notCDom_absSigSum[9:8]; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_5 = |notCDom_absSigSum[11:10]; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_6 = |notCDom_absSigSum[13:12]; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_7 = |notCDom_absSigSum[15:14]; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_8 = |notCDom_absSigSum[17:16]; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_9 = |notCDom_absSigSum[19:18]; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_10 = |notCDom_absSigSum[21:20]; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_11 = |notCDom_absSigSum[23:22]; // @[primitives.scala 104:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_12 = |notCDom_absSigSum[24]; // @[primitives.scala 107:57]
  wire [5:0] notCDom_reduced2AbsSigSum_lo = {notCDom_reduced2AbsSigSum_reducedVec_5,
    notCDom_reduced2AbsSigSum_reducedVec_4,notCDom_reduced2AbsSigSum_reducedVec_3,notCDom_reduced2AbsSigSum_reducedVec_2
    ,notCDom_reduced2AbsSigSum_reducedVec_1,notCDom_reduced2AbsSigSum_reducedVec_0}; // @[primitives.scala 108:20]
  wire [12:0] notCDom_reduced2AbsSigSum = {notCDom_reduced2AbsSigSum_reducedVec_12,
    notCDom_reduced2AbsSigSum_reducedVec_11,notCDom_reduced2AbsSigSum_reducedVec_10,
    notCDom_reduced2AbsSigSum_reducedVec_9,notCDom_reduced2AbsSigSum_reducedVec_8,notCDom_reduced2AbsSigSum_reducedVec_7
    ,notCDom_reduced2AbsSigSum_reducedVec_6,notCDom_reduced2AbsSigSum_lo}; // @[primitives.scala 108:20]
  wire [3:0] _notCDom_normDistReduced2_T_13 = notCDom_reduced2AbsSigSum[1] ? 4'hb : 4'hc; // @[Mux.scala 47:69]
  wire [3:0] _notCDom_normDistReduced2_T_14 = notCDom_reduced2AbsSigSum[2] ? 4'ha : _notCDom_normDistReduced2_T_13; // @[Mux.scala 47:69]
  wire [3:0] _notCDom_normDistReduced2_T_15 = notCDom_reduced2AbsSigSum[3] ? 4'h9 : _notCDom_normDistReduced2_T_14; // @[Mux.scala 47:69]
  wire [3:0] _notCDom_normDistReduced2_T_16 = notCDom_reduced2AbsSigSum[4] ? 4'h8 : _notCDom_normDistReduced2_T_15; // @[Mux.scala 47:69]
  wire [3:0] _notCDom_normDistReduced2_T_17 = notCDom_reduced2AbsSigSum[5] ? 4'h7 : _notCDom_normDistReduced2_T_16; // @[Mux.scala 47:69]
  wire [3:0] _notCDom_normDistReduced2_T_18 = notCDom_reduced2AbsSigSum[6] ? 4'h6 : _notCDom_normDistReduced2_T_17; // @[Mux.scala 47:69]
  wire [3:0] _notCDom_normDistReduced2_T_19 = notCDom_reduced2AbsSigSum[7] ? 4'h5 : _notCDom_normDistReduced2_T_18; // @[Mux.scala 47:69]
  wire [3:0] _notCDom_normDistReduced2_T_20 = notCDom_reduced2AbsSigSum[8] ? 4'h4 : _notCDom_normDistReduced2_T_19; // @[Mux.scala 47:69]
  wire [3:0] _notCDom_normDistReduced2_T_21 = notCDom_reduced2AbsSigSum[9] ? 4'h3 : _notCDom_normDistReduced2_T_20; // @[Mux.scala 47:69]
  wire [3:0] _notCDom_normDistReduced2_T_22 = notCDom_reduced2AbsSigSum[10] ? 4'h2 : _notCDom_normDistReduced2_T_21; // @[Mux.scala 47:69]
  wire [3:0] _notCDom_normDistReduced2_T_23 = notCDom_reduced2AbsSigSum[11] ? 4'h1 : _notCDom_normDistReduced2_T_22; // @[Mux.scala 47:69]
  wire [3:0] notCDom_normDistReduced2 = notCDom_reduced2AbsSigSum[12] ? 4'h0 : _notCDom_normDistReduced2_T_23; // @[Mux.scala 47:69]
  wire [4:0] notCDom_nearNormDist = {notCDom_normDistReduced2, 1'h0}; // @[MulAddRecFN.scala 244:56]
  wire [5:0] _notCDom_sExp_T = {1'b0,$signed(notCDom_nearNormDist)}; // @[MulAddRecFN.scala 245:69]
  wire [6:0] _GEN_4 = {{1{_notCDom_sExp_T[5]}},_notCDom_sExp_T}; // @[MulAddRecFN.scala 245:46]
  wire [6:0] notCDom_sExp = $signed(io_fromPreMul_sExpSum) - $signed(_GEN_4); // @[MulAddRecFN.scala 245:46]
  wire [55:0] _GEN_5 = {{31'd0}, notCDom_absSigSum}; // @[MulAddRecFN.scala 247:27]
  wire [55:0] _notCDom_mainSig_T = _GEN_5 << notCDom_nearNormDist; // @[MulAddRecFN.scala 247:27]
  wire [15:0] notCDom_mainSig = _notCDom_mainSig_T[25:10]; // @[MulAddRecFN.scala 247:50]
  wire [6:0] _notCDom_reduced4SigExtra_T_1 = {notCDom_reduced2AbsSigSum[5:0], 1'h0}; // @[MulAddRecFN.scala 251:55]
  wire  notCDom_reduced4SigExtra_reducedVec_0 = |_notCDom_reduced4SigExtra_T_1[1:0]; // @[primitives.scala 104:54]
  wire  notCDom_reduced4SigExtra_reducedVec_1 = |_notCDom_reduced4SigExtra_T_1[3:2]; // @[primitives.scala 104:54]
  wire  notCDom_reduced4SigExtra_reducedVec_2 = |_notCDom_reduced4SigExtra_T_1[5:4]; // @[primitives.scala 104:54]
  wire  notCDom_reduced4SigExtra_reducedVec_3 = |_notCDom_reduced4SigExtra_T_1[6]; // @[primitives.scala 107:57]
  wire [3:0] _notCDom_reduced4SigExtra_T_2 = {notCDom_reduced4SigExtra_reducedVec_3,
    notCDom_reduced4SigExtra_reducedVec_2,notCDom_reduced4SigExtra_reducedVec_1,notCDom_reduced4SigExtra_reducedVec_0}; // @[primitives.scala 108:20]
  wire [2:0] _notCDom_reduced4SigExtra_T_4 = ~notCDom_normDistReduced2[3:1]; // @[primitives.scala 51:21]
  wire [8:0] notCDom_reduced4SigExtra_shift = 9'sh100 >>> _notCDom_reduced4SigExtra_T_4; // @[primitives.scala 77:58]
  wire  notCDom_reduced4SigExtra_hi_1 = notCDom_reduced4SigExtra_shift[1]; // @[Bitwise.scala 109:18]
  wire  notCDom_reduced4SigExtra_lo_1 = notCDom_reduced4SigExtra_shift[2]; // @[Bitwise.scala 109:44]
  wire  notCDom_reduced4SigExtra_lo_2 = notCDom_reduced4SigExtra_shift[3]; // @[Bitwise.scala 109:44]
  wire [2:0] _notCDom_reduced4SigExtra_T_7 = {notCDom_reduced4SigExtra_hi_1,notCDom_reduced4SigExtra_lo_1,
    notCDom_reduced4SigExtra_lo_2}; // @[Cat.scala 30:58]
  wire [3:0] _GEN_6 = {{1'd0}, _notCDom_reduced4SigExtra_T_7}; // @[MulAddRecFN.scala 251:78]
  wire [3:0] _notCDom_reduced4SigExtra_T_8 = _notCDom_reduced4SigExtra_T_2 & _GEN_6; // @[MulAddRecFN.scala 251:78]
  wire  notCDom_reduced4SigExtra = |_notCDom_reduced4SigExtra_T_8; // @[MulAddRecFN.scala 253:11]
  wire [12:0] notCDom_sig_hi = notCDom_mainSig[15:3]; // @[MulAddRecFN.scala 255:28]
  wire  notCDom_sig_lo = |notCDom_mainSig[2:0] | notCDom_reduced4SigExtra; // @[MulAddRecFN.scala 256:39]
  wire [13:0] notCDom_sig = {notCDom_sig_hi,notCDom_sig_lo}; // @[Cat.scala 30:58]
  wire  notCDom_completeCancellation = notCDom_sig[13:12] == 2'h0; // @[MulAddRecFN.scala 259:50]
  wire  _notCDom_sign_T = io_fromPreMul_signProd ^ notCDom_signSigSum; // @[MulAddRecFN.scala 263:36]
  wire  notCDom_sign = notCDom_completeCancellation ? 1'h0 : _notCDom_sign_T; // @[MulAddRecFN.scala 261:12]
  wire  notNaN_isInfProd = io_fromPreMul_isInfA | io_fromPreMul_isInfB; // @[MulAddRecFN.scala 268:49]
  wire  notNaN_isInfOut = notNaN_isInfProd | io_fromPreMul_isInfC; // @[MulAddRecFN.scala 269:44]
  wire  notNaN_addZeros = (io_fromPreMul_isZeroA | io_fromPreMul_isZeroB) & io_fromPreMul_isZeroC; // @[MulAddRecFN.scala 271:58]
  wire  _io_invalidExc_T = io_fromPreMul_isInfA & io_fromPreMul_isZeroB; // @[MulAddRecFN.scala 276:31]
  wire  _io_invalidExc_T_1 = io_fromPreMul_isSigNaNAny | _io_invalidExc_T; // @[MulAddRecFN.scala 275:35]
  wire  _io_invalidExc_T_2 = io_fromPreMul_isZeroA & io_fromPreMul_isInfB; // @[MulAddRecFN.scala 277:32]
  wire  _io_invalidExc_T_3 = _io_invalidExc_T_1 | _io_invalidExc_T_2; // @[MulAddRecFN.scala 276:57]
  wire  _io_invalidExc_T_6 = ~io_fromPreMul_isNaNAOrB & notNaN_isInfProd; // @[MulAddRecFN.scala 278:36]
  wire  _io_invalidExc_T_7 = _io_invalidExc_T_6 & io_fromPreMul_isInfC; // @[MulAddRecFN.scala 279:61]
  wire  _io_invalidExc_T_8 = _io_invalidExc_T_7 & io_fromPreMul_doSubMags; // @[MulAddRecFN.scala 280:35]
  wire  _io_rawOut_isZero_T_1 = ~io_fromPreMul_CIsDominant & notCDom_completeCancellation; // @[MulAddRecFN.scala 287:42]
  wire  _io_rawOut_sign_T_1 = io_fromPreMul_isInfC & CDom_sign; // @[MulAddRecFN.scala 290:31]
  wire  _io_rawOut_sign_T_2 = notNaN_isInfProd & io_fromPreMul_signProd | _io_rawOut_sign_T_1; // @[MulAddRecFN.scala 289:54]
  wire  _io_rawOut_sign_T_5 = notNaN_addZeros & io_fromPreMul_signProd; // @[MulAddRecFN.scala 291:48]
  wire  _io_rawOut_sign_T_6 = _io_rawOut_sign_T_5 & CDom_sign; // @[MulAddRecFN.scala 292:36]
  wire  _io_rawOut_sign_T_7 = _io_rawOut_sign_T_2 | _io_rawOut_sign_T_6; // @[MulAddRecFN.scala 290:43]
  wire  _io_rawOut_sign_T_15 = io_fromPreMul_CIsDominant ? CDom_sign : notCDom_sign; // @[MulAddRecFN.scala 296:17]
  wire  _io_rawOut_sign_T_16 = ~notNaN_isInfOut & ~notNaN_addZeros & _io_rawOut_sign_T_15; // @[MulAddRecFN.scala 295:49]
  assign io_invalidExc = _io_invalidExc_T_3 | _io_invalidExc_T_8; // @[MulAddRecFN.scala 277:57]
  assign io_rawOut_isNaN = io_fromPreMul_isNaNAOrB | io_fromPreMul_isNaNC; // @[MulAddRecFN.scala 282:48]
  assign io_rawOut_isInf = notNaN_isInfProd | io_fromPreMul_isInfC; // @[MulAddRecFN.scala 269:44]
  assign io_rawOut_isZero = notNaN_addZeros | _io_rawOut_isZero_T_1; // @[MulAddRecFN.scala 286:25]
  assign io_rawOut_sign = _io_rawOut_sign_T_7 | _io_rawOut_sign_T_16; // @[MulAddRecFN.scala 294:50]
  assign io_rawOut_sExp = io_fromPreMul_CIsDominant ? $signed(CDom_sExp) : $signed(notCDom_sExp); // @[MulAddRecFN.scala 297:26]
  assign io_rawOut_sig = io_fromPreMul_CIsDominant ? CDom_sig : notCDom_sig; // @[MulAddRecFN.scala 298:25]
endmodule
module RoundAnyRawFNToRecFN(
  input         io_invalidExc,
  input         io_in_isNaN,
  input         io_in_isInf,
  input         io_in_isZero,
  input         io_in_sign,
  input  [6:0]  io_in_sExp,
  input  [13:0] io_in_sig,
  output [16:0] io_out
);
  wire  doShiftSigDown1 = io_in_sig[13]; // @[RoundAnyRawFNToRecFN.scala 118:61]
  wire [5:0] _roundMask_T_1 = ~io_in_sExp[5:0]; // @[primitives.scala 51:21]
  wire [64:0] roundMask_shift = 65'sh10000000000000000 >>> _roundMask_T_1; // @[primitives.scala 77:58]
  wire [7:0] _roundMask_T_7 = {{4'd0}, roundMask_shift[14:11]}; // @[Bitwise.scala 103:31]
  wire [7:0] _roundMask_T_9 = {roundMask_shift[10:7], 4'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _roundMask_T_11 = _roundMask_T_9 & 8'hf0; // @[Bitwise.scala 103:75]
  wire [7:0] _roundMask_T_12 = _roundMask_T_7 | _roundMask_T_11; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_0 = {{2'd0}, _roundMask_T_12[7:2]}; // @[Bitwise.scala 103:31]
  wire [7:0] _roundMask_T_17 = _GEN_0 & 8'h33; // @[Bitwise.scala 103:31]
  wire [7:0] _roundMask_T_19 = {_roundMask_T_12[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _roundMask_T_21 = _roundMask_T_19 & 8'hcc; // @[Bitwise.scala 103:75]
  wire [7:0] _roundMask_T_22 = _roundMask_T_17 | _roundMask_T_21; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_1 = {{1'd0}, _roundMask_T_22[7:1]}; // @[Bitwise.scala 103:31]
  wire [7:0] _roundMask_T_27 = _GEN_1 & 8'h55; // @[Bitwise.scala 103:31]
  wire [7:0] _roundMask_T_29 = {_roundMask_T_22[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _roundMask_T_31 = _roundMask_T_29 & 8'haa; // @[Bitwise.scala 103:75]
  wire [7:0] roundMask_hi = _roundMask_T_27 | _roundMask_T_31; // @[Bitwise.scala 103:39]
  wire  roundMask_hi_1 = roundMask_shift[15]; // @[Bitwise.scala 109:18]
  wire  roundMask_lo = roundMask_shift[16]; // @[Bitwise.scala 109:44]
  wire  roundMask_hi_3 = roundMask_shift[17]; // @[Bitwise.scala 109:18]
  wire  roundMask_lo_1 = roundMask_shift[18]; // @[Bitwise.scala 109:44]
  wire [11:0] _roundMask_T_35 = {roundMask_hi,roundMask_hi_1,roundMask_lo,roundMask_hi_3,roundMask_lo_1}; // @[Cat.scala 30:58]
  wire [11:0] _GEN_2 = {{11'd0}, doShiftSigDown1}; // @[RoundAnyRawFNToRecFN.scala 157:23]
  wire [11:0] roundMask_hi_4 = _roundMask_T_35 | _GEN_2; // @[RoundAnyRawFNToRecFN.scala 157:23]
  wire [13:0] roundMask = {roundMask_hi_4,2'h3}; // @[Cat.scala 30:58]
  wire [12:0] shiftedRoundMask_lo = roundMask[13:1]; // @[RoundAnyRawFNToRecFN.scala 160:57]
  wire [13:0] shiftedRoundMask = {1'h0,shiftedRoundMask_lo}; // @[Cat.scala 30:58]
  wire [13:0] _roundPosMask_T = ~shiftedRoundMask; // @[RoundAnyRawFNToRecFN.scala 161:28]
  wire [13:0] roundPosMask = _roundPosMask_T & roundMask; // @[RoundAnyRawFNToRecFN.scala 161:46]
  wire [13:0] _roundPosBit_T = io_in_sig & roundPosMask; // @[RoundAnyRawFNToRecFN.scala 162:40]
  wire  roundPosBit = |_roundPosBit_T; // @[RoundAnyRawFNToRecFN.scala 162:56]
  wire [13:0] _anyRoundExtra_T = io_in_sig & shiftedRoundMask; // @[RoundAnyRawFNToRecFN.scala 163:42]
  wire  anyRoundExtra = |_anyRoundExtra_T; // @[RoundAnyRawFNToRecFN.scala 163:62]
  wire [13:0] _roundedSig_T = io_in_sig | roundMask; // @[RoundAnyRawFNToRecFN.scala 172:32]
  wire [12:0] _roundedSig_T_2 = _roundedSig_T[13:2] + 12'h1; // @[RoundAnyRawFNToRecFN.scala 172:49]
  wire  _roundedSig_T_4 = ~anyRoundExtra; // @[RoundAnyRawFNToRecFN.scala 174:30]
  wire [12:0] _roundedSig_T_7 = roundPosBit & _roundedSig_T_4 ? shiftedRoundMask_lo : 13'h0; // @[RoundAnyRawFNToRecFN.scala 173:25]
  wire [12:0] _roundedSig_T_8 = ~_roundedSig_T_7; // @[RoundAnyRawFNToRecFN.scala 173:21]
  wire [12:0] _roundedSig_T_9 = _roundedSig_T_2 & _roundedSig_T_8; // @[RoundAnyRawFNToRecFN.scala 172:61]
  wire [13:0] _roundedSig_T_10 = ~roundMask; // @[RoundAnyRawFNToRecFN.scala 178:32]
  wire [13:0] _roundedSig_T_11 = io_in_sig & _roundedSig_T_10; // @[RoundAnyRawFNToRecFN.scala 178:30]
  wire [12:0] _roundedSig_T_16 = {{1'd0}, _roundedSig_T_11[13:2]}; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [12:0] roundedSig = roundPosBit ? _roundedSig_T_9 : _roundedSig_T_16; // @[RoundAnyRawFNToRecFN.scala 171:16]
  wire [2:0] _sRoundedExp_T_1 = {1'b0,$signed(roundedSig[12:11])}; // @[RoundAnyRawFNToRecFN.scala 183:69]
  wire [6:0] _GEN_3 = {{4{_sRoundedExp_T_1[2]}},_sRoundedExp_T_1}; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [7:0] sRoundedExp = $signed(io_in_sExp) + $signed(_GEN_3); // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [5:0] common_expOut = sRoundedExp[5:0]; // @[RoundAnyRawFNToRecFN.scala 185:37]
  wire [9:0] common_fractOut = doShiftSigDown1 ? roundedSig[10:1] : roundedSig[9:0]; // @[RoundAnyRawFNToRecFN.scala 187:16]
  wire [3:0] _common_overflow_T = sRoundedExp[7:4]; // @[RoundAnyRawFNToRecFN.scala 194:30]
  wire  common_overflow = $signed(_common_overflow_T) >= 4'sh3; // @[RoundAnyRawFNToRecFN.scala 194:50]
  wire  common_totalUnderflow = $signed(sRoundedExp) < 8'sh8; // @[RoundAnyRawFNToRecFN.scala 198:31]
  wire  isNaNOut = io_invalidExc | io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 233:34]
  wire  commonCase = ~isNaNOut & ~io_in_isInf & ~io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 235:61]
  wire  overflow = commonCase & common_overflow; // @[RoundAnyRawFNToRecFN.scala 236:32]
  wire  notNaN_isInfOut = io_in_isInf | overflow; // @[RoundAnyRawFNToRecFN.scala 246:32]
  wire  signOut = isNaNOut ? 1'h0 : io_in_sign; // @[RoundAnyRawFNToRecFN.scala 248:22]
  wire [5:0] _expOut_T_1 = io_in_isZero | common_totalUnderflow ? 6'h38 : 6'h0; // @[RoundAnyRawFNToRecFN.scala 251:18]
  wire [5:0] _expOut_T_2 = ~_expOut_T_1; // @[RoundAnyRawFNToRecFN.scala 251:14]
  wire [5:0] _expOut_T_3 = common_expOut & _expOut_T_2; // @[RoundAnyRawFNToRecFN.scala 250:24]
  wire [5:0] _expOut_T_11 = notNaN_isInfOut ? 6'h8 : 6'h0; // @[RoundAnyRawFNToRecFN.scala 263:18]
  wire [5:0] _expOut_T_12 = ~_expOut_T_11; // @[RoundAnyRawFNToRecFN.scala 263:14]
  wire [5:0] _expOut_T_13 = _expOut_T_3 & _expOut_T_12; // @[RoundAnyRawFNToRecFN.scala 262:17]
  wire [5:0] _expOut_T_18 = notNaN_isInfOut ? 6'h30 : 6'h0; // @[RoundAnyRawFNToRecFN.scala 275:16]
  wire [5:0] _expOut_T_19 = _expOut_T_13 | _expOut_T_18; // @[RoundAnyRawFNToRecFN.scala 274:15]
  wire [5:0] _expOut_T_20 = isNaNOut ? 6'h38 : 6'h0; // @[RoundAnyRawFNToRecFN.scala 276:16]
  wire [5:0] expOut = _expOut_T_19 | _expOut_T_20; // @[RoundAnyRawFNToRecFN.scala 275:77]
  wire [9:0] _fractOut_T_2 = isNaNOut ? 10'h200 : 10'h0; // @[RoundAnyRawFNToRecFN.scala 279:16]
  wire [9:0] fractOut = isNaNOut | io_in_isZero | common_totalUnderflow ? _fractOut_T_2 : common_fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12]
  wire [6:0] io_out_hi = {signOut,expOut}; // @[Cat.scala 30:58]
  assign io_out = {io_out_hi,fractOut}; // @[Cat.scala 30:58]
endmodule
module RoundRawFNToRecFN(
  input         io_invalidExc,
  input         io_in_isNaN,
  input         io_in_isInf,
  input         io_in_isZero,
  input         io_in_sign,
  input  [6:0]  io_in_sExp,
  input  [13:0] io_in_sig,
  output [16:0] io_out
);
  wire  roundAnyRawFNToRecFN_io_invalidExc; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_sign; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [6:0] roundAnyRawFNToRecFN_io_in_sExp; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [13:0] roundAnyRawFNToRecFN_io_in_sig; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [16:0] roundAnyRawFNToRecFN_io_out; // @[RoundAnyRawFNToRecFN.scala 307:15]
  RoundAnyRawFNToRecFN roundAnyRawFNToRecFN ( // @[RoundAnyRawFNToRecFN.scala 307:15]
    .io_invalidExc(roundAnyRawFNToRecFN_io_invalidExc),
    .io_in_isNaN(roundAnyRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundAnyRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundAnyRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundAnyRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundAnyRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundAnyRawFNToRecFN_io_in_sig),
    .io_out(roundAnyRawFNToRecFN_io_out)
  );
  assign io_out = roundAnyRawFNToRecFN_io_out; // @[RoundAnyRawFNToRecFN.scala 315:23]
  assign roundAnyRawFNToRecFN_io_invalidExc = io_invalidExc; // @[RoundAnyRawFNToRecFN.scala 310:44]
  assign roundAnyRawFNToRecFN_io_in_isNaN = io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_isInf = io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_isZero = io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_sign = io_in_sign; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_sExp = io_in_sExp; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_sig = io_in_sig; // @[RoundAnyRawFNToRecFN.scala 312:44]
endmodule
module MulAddRecFN(
  input  [16:0] io_a,
  input  [16:0] io_b,
  input  [16:0] io_c,
  output [16:0] io_out,
  output [21:0] io_mulOut,
  output [21:0] io_mulIn1,
  output [21:0] io_mulIn2,
  output        io_correctMulOut,
  output        io_correctMulIn,
  output        io_sigSum_Msb
);
  wire [16:0] mulAddRecFNToRaw_preMul_io_a; // @[MulAddRecFN.scala 327:15]
  wire [16:0] mulAddRecFNToRaw_preMul_io_b; // @[MulAddRecFN.scala 327:15]
  wire [16:0] mulAddRecFNToRaw_preMul_io_c; // @[MulAddRecFN.scala 327:15]
  wire [10:0] mulAddRecFNToRaw_preMul_io_mulAddA; // @[MulAddRecFN.scala 327:15]
  wire [10:0] mulAddRecFNToRaw_preMul_io_mulAddB; // @[MulAddRecFN.scala 327:15]
  wire [21:0] mulAddRecFNToRaw_preMul_io_mulAddC; // @[MulAddRecFN.scala 327:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny; // @[MulAddRecFN.scala 327:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB; // @[MulAddRecFN.scala 327:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfA; // @[MulAddRecFN.scala 327:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA; // @[MulAddRecFN.scala 327:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfB; // @[MulAddRecFN.scala 327:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB; // @[MulAddRecFN.scala 327:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_signProd; // @[MulAddRecFN.scala 327:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC; // @[MulAddRecFN.scala 327:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfC; // @[MulAddRecFN.scala 327:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC; // @[MulAddRecFN.scala 327:15]
  wire [6:0] mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum; // @[MulAddRecFN.scala 327:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags; // @[MulAddRecFN.scala 327:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant; // @[MulAddRecFN.scala 327:15]
  wire [3:0] mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist; // @[MulAddRecFN.scala 327:15]
  wire [12:0] mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC; // @[MulAddRecFN.scala 327:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC; // @[MulAddRecFN.scala 327:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny; // @[MulAddRecFN.scala 329:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB; // @[MulAddRecFN.scala 329:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA; // @[MulAddRecFN.scala 329:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA; // @[MulAddRecFN.scala 329:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB; // @[MulAddRecFN.scala 329:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB; // @[MulAddRecFN.scala 329:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_signProd; // @[MulAddRecFN.scala 329:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC; // @[MulAddRecFN.scala 329:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC; // @[MulAddRecFN.scala 329:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC; // @[MulAddRecFN.scala 329:15]
  wire [6:0] mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum; // @[MulAddRecFN.scala 329:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags; // @[MulAddRecFN.scala 329:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant; // @[MulAddRecFN.scala 329:15]
  wire [3:0] mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist; // @[MulAddRecFN.scala 329:15]
  wire [12:0] mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC; // @[MulAddRecFN.scala 329:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC; // @[MulAddRecFN.scala 329:15]
  wire [22:0] mulAddRecFNToRaw_postMul_io_mulAddResult; // @[MulAddRecFN.scala 329:15]
  wire  mulAddRecFNToRaw_postMul_io_invalidExc; // @[MulAddRecFN.scala 329:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isNaN; // @[MulAddRecFN.scala 329:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isInf; // @[MulAddRecFN.scala 329:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isZero; // @[MulAddRecFN.scala 329:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_sign; // @[MulAddRecFN.scala 329:15]
  wire [6:0] mulAddRecFNToRaw_postMul_io_rawOut_sExp; // @[MulAddRecFN.scala 329:15]
  wire [13:0] mulAddRecFNToRaw_postMul_io_rawOut_sig; // @[MulAddRecFN.scala 329:15]
  wire  roundRawFNToRecFN_io_invalidExc; // @[MulAddRecFN.scala 369:15]
  wire  roundRawFNToRecFN_io_in_isNaN; // @[MulAddRecFN.scala 369:15]
  wire  roundRawFNToRecFN_io_in_isInf; // @[MulAddRecFN.scala 369:15]
  wire  roundRawFNToRecFN_io_in_isZero; // @[MulAddRecFN.scala 369:15]
  wire  roundRawFNToRecFN_io_in_sign; // @[MulAddRecFN.scala 369:15]
  wire [6:0] roundRawFNToRecFN_io_in_sExp; // @[MulAddRecFN.scala 369:15]
  wire [13:0] roundRawFNToRecFN_io_in_sig; // @[MulAddRecFN.scala 369:15]
  wire [16:0] roundRawFNToRecFN_io_out; // @[MulAddRecFN.scala 369:15]
  wire  _io_correctMulOut_T_1 = io_mulOut >= 22'h100000; // @[MulAddRecFN.scala 344:17]
  wire [22:0] mulAddResult = io_mulOut + mulAddRecFNToRaw_preMul_io_mulAddC; // @[MulAddRecFN.scala 350:21]
  MulAddRecFNToRaw_preMul mulAddRecFNToRaw_preMul ( // @[MulAddRecFN.scala 327:15]
    .io_a(mulAddRecFNToRaw_preMul_io_a),
    .io_b(mulAddRecFNToRaw_preMul_io_b),
    .io_c(mulAddRecFNToRaw_preMul_io_c),
    .io_mulAddA(mulAddRecFNToRaw_preMul_io_mulAddA),
    .io_mulAddB(mulAddRecFNToRaw_preMul_io_mulAddB),
    .io_mulAddC(mulAddRecFNToRaw_preMul_io_mulAddC),
    .io_toPostMul_isSigNaNAny(mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny),
    .io_toPostMul_isNaNAOrB(mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB),
    .io_toPostMul_isInfA(mulAddRecFNToRaw_preMul_io_toPostMul_isInfA),
    .io_toPostMul_isZeroA(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA),
    .io_toPostMul_isInfB(mulAddRecFNToRaw_preMul_io_toPostMul_isInfB),
    .io_toPostMul_isZeroB(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB),
    .io_toPostMul_signProd(mulAddRecFNToRaw_preMul_io_toPostMul_signProd),
    .io_toPostMul_isNaNC(mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC),
    .io_toPostMul_isInfC(mulAddRecFNToRaw_preMul_io_toPostMul_isInfC),
    .io_toPostMul_isZeroC(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC),
    .io_toPostMul_sExpSum(mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum),
    .io_toPostMul_doSubMags(mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags),
    .io_toPostMul_CIsDominant(mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant),
    .io_toPostMul_CDom_CAlignDist(mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist),
    .io_toPostMul_highAlignedSigC(mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC),
    .io_toPostMul_bit0AlignedSigC(mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC)
  );
  MulAddRecFNToRaw_postMul mulAddRecFNToRaw_postMul ( // @[MulAddRecFN.scala 329:15]
    .io_fromPreMul_isSigNaNAny(mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny),
    .io_fromPreMul_isNaNAOrB(mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB),
    .io_fromPreMul_isInfA(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA),
    .io_fromPreMul_isZeroA(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA),
    .io_fromPreMul_isInfB(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB),
    .io_fromPreMul_isZeroB(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB),
    .io_fromPreMul_signProd(mulAddRecFNToRaw_postMul_io_fromPreMul_signProd),
    .io_fromPreMul_isNaNC(mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC),
    .io_fromPreMul_isInfC(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC),
    .io_fromPreMul_isZeroC(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC),
    .io_fromPreMul_sExpSum(mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum),
    .io_fromPreMul_doSubMags(mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags),
    .io_fromPreMul_CIsDominant(mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant),
    .io_fromPreMul_CDom_CAlignDist(mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist),
    .io_fromPreMul_highAlignedSigC(mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC),
    .io_fromPreMul_bit0AlignedSigC(mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC),
    .io_mulAddResult(mulAddRecFNToRaw_postMul_io_mulAddResult),
    .io_invalidExc(mulAddRecFNToRaw_postMul_io_invalidExc),
    .io_rawOut_isNaN(mulAddRecFNToRaw_postMul_io_rawOut_isNaN),
    .io_rawOut_isInf(mulAddRecFNToRaw_postMul_io_rawOut_isInf),
    .io_rawOut_isZero(mulAddRecFNToRaw_postMul_io_rawOut_isZero),
    .io_rawOut_sign(mulAddRecFNToRaw_postMul_io_rawOut_sign),
    .io_rawOut_sExp(mulAddRecFNToRaw_postMul_io_rawOut_sExp),
    .io_rawOut_sig(mulAddRecFNToRaw_postMul_io_rawOut_sig)
  );
  RoundRawFNToRecFN roundRawFNToRecFN ( // @[MulAddRecFN.scala 369:15]
    .io_invalidExc(roundRawFNToRecFN_io_invalidExc),
    .io_in_isNaN(roundRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundRawFNToRecFN_io_in_sig),
    .io_out(roundRawFNToRecFN_io_out)
  );
  assign io_out = roundRawFNToRecFN_io_out; // @[MulAddRecFN.scala 375:23]
  assign io_mulOut = mulAddRecFNToRaw_preMul_io_mulAddA * mulAddRecFNToRaw_preMul_io_mulAddB; // @[MulAddRecFN.scala 336:54]
  assign io_mulIn1 = {{11'd0}, mulAddRecFNToRaw_preMul_io_mulAddA}; // @[MulAddRecFN.scala 339:15]
  assign io_mulIn2 = {{11'd0}, mulAddRecFNToRaw_preMul_io_mulAddB}; // @[MulAddRecFN.scala 340:15]
  assign io_correctMulOut = io_mulOut <= 22'h3ff001 & _io_correctMulOut_T_1; // @[MulAddRecFN.scala 343:84]
  assign io_correctMulIn = io_mulIn1[10] & io_mulIn2[10]; // @[MulAddRecFN.scala 347:41]
  assign io_sigSum_Msb = mulAddResult[22]; // @[MulAddRecFN.scala 353:34]
  assign mulAddRecFNToRaw_preMul_io_a = io_a; // @[MulAddRecFN.scala 332:35]
  assign mulAddRecFNToRaw_preMul_io_b = io_b; // @[MulAddRecFN.scala 333:35]
  assign mulAddRecFNToRaw_preMul_io_c = io_c; // @[MulAddRecFN.scala 334:35]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny = mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny; // @[MulAddRecFN.scala 361:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB = mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB; // @[MulAddRecFN.scala 361:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA = mulAddRecFNToRaw_preMul_io_toPostMul_isInfA; // @[MulAddRecFN.scala 361:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA = mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA; // @[MulAddRecFN.scala 361:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB = mulAddRecFNToRaw_preMul_io_toPostMul_isInfB; // @[MulAddRecFN.scala 361:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB = mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB; // @[MulAddRecFN.scala 361:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_signProd = mulAddRecFNToRaw_preMul_io_toPostMul_signProd; // @[MulAddRecFN.scala 361:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC = mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC; // @[MulAddRecFN.scala 361:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC = mulAddRecFNToRaw_preMul_io_toPostMul_isInfC; // @[MulAddRecFN.scala 361:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC = mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC; // @[MulAddRecFN.scala 361:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum = mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum; // @[MulAddRecFN.scala 361:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags = mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags; // @[MulAddRecFN.scala 361:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant = mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant; // @[MulAddRecFN.scala 361:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist = mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist; // @[MulAddRecFN.scala 361:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC = mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC; // @[MulAddRecFN.scala 361:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC = mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC; // @[MulAddRecFN.scala 361:44]
  assign mulAddRecFNToRaw_postMul_io_mulAddResult = io_mulOut + mulAddRecFNToRaw_preMul_io_mulAddC; // @[MulAddRecFN.scala 350:21]
  assign roundRawFNToRecFN_io_invalidExc = mulAddRecFNToRaw_postMul_io_invalidExc; // @[MulAddRecFN.scala 370:39]
  assign roundRawFNToRecFN_io_in_isNaN = mulAddRecFNToRaw_postMul_io_rawOut_isNaN; // @[MulAddRecFN.scala 372:39]
  assign roundRawFNToRecFN_io_in_isInf = mulAddRecFNToRaw_postMul_io_rawOut_isInf; // @[MulAddRecFN.scala 372:39]
  assign roundRawFNToRecFN_io_in_isZero = mulAddRecFNToRaw_postMul_io_rawOut_isZero; // @[MulAddRecFN.scala 372:39]
  assign roundRawFNToRecFN_io_in_sign = mulAddRecFNToRaw_postMul_io_rawOut_sign; // @[MulAddRecFN.scala 372:39]
  assign roundRawFNToRecFN_io_in_sExp = mulAddRecFNToRaw_postMul_io_rawOut_sExp; // @[MulAddRecFN.scala 372:39]
  assign roundRawFNToRecFN_io_in_sig = mulAddRecFNToRaw_postMul_io_rawOut_sig; // @[MulAddRecFN.scala 372:39]
endmodule
module FP16MulAdder(
  input  [15:0] io_a,
  input  [15:0] io_b,
  input  [15:0] io_c,
  output [15:0] io_out
);
  wire [16:0] mulAddRecFN_io_a; // @[hardfloat.scala 31:29]
  wire [16:0] mulAddRecFN_io_b; // @[hardfloat.scala 31:29]
  wire [16:0] mulAddRecFN_io_c; // @[hardfloat.scala 31:29]
  wire [16:0] mulAddRecFN_io_out; // @[hardfloat.scala 31:29]
  wire [21:0] mulAddRecFN_io_mulOut; // @[hardfloat.scala 31:29]
  wire [21:0] mulAddRecFN_io_mulIn1; // @[hardfloat.scala 31:29]
  wire [21:0] mulAddRecFN_io_mulIn2; // @[hardfloat.scala 31:29]
  wire  mulAddRecFN_io_correctMulOut; // @[hardfloat.scala 31:29]
  wire  mulAddRecFN_io_correctMulIn; // @[hardfloat.scala 31:29]
  wire  mulAddRecFN_io_sigSum_Msb; // @[hardfloat.scala 31:29]
  wire  mulAddRecFN_io_a_rawIn_sign = io_a[15]; // @[rawFloatFromFN.scala 46:22]
  wire [4:0] mulAddRecFN_io_a_rawIn_expIn = io_a[14:10]; // @[rawFloatFromFN.scala 47:23]
  wire [9:0] mulAddRecFN_io_a_rawIn_fractIn = io_a[9:0]; // @[rawFloatFromFN.scala 48:25]
  wire  mulAddRecFN_io_a_rawIn_isZeroExpIn = mulAddRecFN_io_a_rawIn_expIn == 5'h0; // @[rawFloatFromFN.scala 50:34]
  wire  mulAddRecFN_io_a_rawIn_isZeroFractIn = mulAddRecFN_io_a_rawIn_fractIn == 10'h0; // @[rawFloatFromFN.scala 51:38]
  wire [3:0] _mulAddRecFN_io_a_rawIn_normDist_T_10 = mulAddRecFN_io_a_rawIn_fractIn[1] ? 4'h8 : 4'h9; // @[Mux.scala 47:69]
  wire [3:0] _mulAddRecFN_io_a_rawIn_normDist_T_11 = mulAddRecFN_io_a_rawIn_fractIn[2] ? 4'h7 :
    _mulAddRecFN_io_a_rawIn_normDist_T_10; // @[Mux.scala 47:69]
  wire [3:0] _mulAddRecFN_io_a_rawIn_normDist_T_12 = mulAddRecFN_io_a_rawIn_fractIn[3] ? 4'h6 :
    _mulAddRecFN_io_a_rawIn_normDist_T_11; // @[Mux.scala 47:69]
  wire [3:0] _mulAddRecFN_io_a_rawIn_normDist_T_13 = mulAddRecFN_io_a_rawIn_fractIn[4] ? 4'h5 :
    _mulAddRecFN_io_a_rawIn_normDist_T_12; // @[Mux.scala 47:69]
  wire [3:0] _mulAddRecFN_io_a_rawIn_normDist_T_14 = mulAddRecFN_io_a_rawIn_fractIn[5] ? 4'h4 :
    _mulAddRecFN_io_a_rawIn_normDist_T_13; // @[Mux.scala 47:69]
  wire [3:0] _mulAddRecFN_io_a_rawIn_normDist_T_15 = mulAddRecFN_io_a_rawIn_fractIn[6] ? 4'h3 :
    _mulAddRecFN_io_a_rawIn_normDist_T_14; // @[Mux.scala 47:69]
  wire [3:0] _mulAddRecFN_io_a_rawIn_normDist_T_16 = mulAddRecFN_io_a_rawIn_fractIn[7] ? 4'h2 :
    _mulAddRecFN_io_a_rawIn_normDist_T_15; // @[Mux.scala 47:69]
  wire [3:0] _mulAddRecFN_io_a_rawIn_normDist_T_17 = mulAddRecFN_io_a_rawIn_fractIn[8] ? 4'h1 :
    _mulAddRecFN_io_a_rawIn_normDist_T_16; // @[Mux.scala 47:69]
  wire [3:0] mulAddRecFN_io_a_rawIn_normDist = mulAddRecFN_io_a_rawIn_fractIn[9] ? 4'h0 :
    _mulAddRecFN_io_a_rawIn_normDist_T_17; // @[Mux.scala 47:69]
  wire [24:0] _GEN_0 = {{15'd0}, mulAddRecFN_io_a_rawIn_fractIn}; // @[rawFloatFromFN.scala 54:36]
  wire [24:0] _mulAddRecFN_io_a_rawIn_subnormFract_T = _GEN_0 << mulAddRecFN_io_a_rawIn_normDist; // @[rawFloatFromFN.scala 54:36]
  wire [9:0] mulAddRecFN_io_a_rawIn_subnormFract = {_mulAddRecFN_io_a_rawIn_subnormFract_T[8:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  wire [5:0] _GEN_1 = {{2'd0}, mulAddRecFN_io_a_rawIn_normDist}; // @[rawFloatFromFN.scala 57:26]
  wire [5:0] _mulAddRecFN_io_a_rawIn_adjustedExp_T = _GEN_1 ^ 6'h3f; // @[rawFloatFromFN.scala 57:26]
  wire [5:0] _mulAddRecFN_io_a_rawIn_adjustedExp_T_1 = mulAddRecFN_io_a_rawIn_isZeroExpIn ?
    _mulAddRecFN_io_a_rawIn_adjustedExp_T : {{1'd0}, mulAddRecFN_io_a_rawIn_expIn}; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _mulAddRecFN_io_a_rawIn_adjustedExp_T_2 = mulAddRecFN_io_a_rawIn_isZeroExpIn ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  wire [4:0] _GEN_2 = {{3'd0}, _mulAddRecFN_io_a_rawIn_adjustedExp_T_2}; // @[rawFloatFromFN.scala 60:22]
  wire [4:0] _mulAddRecFN_io_a_rawIn_adjustedExp_T_3 = 5'h10 | _GEN_2; // @[rawFloatFromFN.scala 60:22]
  wire [5:0] _GEN_3 = {{1'd0}, _mulAddRecFN_io_a_rawIn_adjustedExp_T_3}; // @[rawFloatFromFN.scala 59:15]
  wire [5:0] mulAddRecFN_io_a_rawIn_adjustedExp = _mulAddRecFN_io_a_rawIn_adjustedExp_T_1 + _GEN_3; // @[rawFloatFromFN.scala 59:15]
  wire  mulAddRecFN_io_a_rawIn_isZero = mulAddRecFN_io_a_rawIn_isZeroExpIn & mulAddRecFN_io_a_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 62:34]
  wire  mulAddRecFN_io_a_rawIn_isSpecial = mulAddRecFN_io_a_rawIn_adjustedExp[5:4] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  wire  mulAddRecFN_io_a_rawIn__isNaN = mulAddRecFN_io_a_rawIn_isSpecial & ~mulAddRecFN_io_a_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 66:33]
  wire [6:0] mulAddRecFN_io_a_rawIn__sExp = {1'b0,$signed(mulAddRecFN_io_a_rawIn_adjustedExp)}; // @[rawFloatFromFN.scala 70:48]
  wire  mulAddRecFN_io_a_rawIn_out_sig_hi_lo = ~mulAddRecFN_io_a_rawIn_isZero; // @[rawFloatFromFN.scala 72:29]
  wire [9:0] mulAddRecFN_io_a_rawIn_out_sig_lo = mulAddRecFN_io_a_rawIn_isZeroExpIn ?
    mulAddRecFN_io_a_rawIn_subnormFract : mulAddRecFN_io_a_rawIn_fractIn; // @[rawFloatFromFN.scala 72:42]
  wire [11:0] mulAddRecFN_io_a_rawIn__sig = {1'h0,mulAddRecFN_io_a_rawIn_out_sig_hi_lo,mulAddRecFN_io_a_rawIn_out_sig_lo
    }; // @[Cat.scala 30:58]
  wire [2:0] _mulAddRecFN_io_a_T_1 = mulAddRecFN_io_a_rawIn_isZero ? 3'h0 : mulAddRecFN_io_a_rawIn__sExp[5:3]; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_4 = {{2'd0}, mulAddRecFN_io_a_rawIn__isNaN}; // @[recFNFromFN.scala 48:79]
  wire [2:0] mulAddRecFN_io_a_hi_lo = _mulAddRecFN_io_a_T_1 | _GEN_4; // @[recFNFromFN.scala 48:79]
  wire [2:0] mulAddRecFN_io_a_lo_hi = mulAddRecFN_io_a_rawIn__sExp[2:0]; // @[recFNFromFN.scala 50:23]
  wire [9:0] mulAddRecFN_io_a_lo_lo = mulAddRecFN_io_a_rawIn__sig[9:0]; // @[recFNFromFN.scala 51:22]
  wire [12:0] mulAddRecFN_io_a_lo = {mulAddRecFN_io_a_lo_hi,mulAddRecFN_io_a_lo_lo}; // @[Cat.scala 30:58]
  wire [3:0] mulAddRecFN_io_a_hi = {mulAddRecFN_io_a_rawIn_sign,mulAddRecFN_io_a_hi_lo}; // @[Cat.scala 30:58]
  wire  mulAddRecFN_io_b_rawIn_sign = io_b[15]; // @[rawFloatFromFN.scala 46:22]
  wire [4:0] mulAddRecFN_io_b_rawIn_expIn = io_b[14:10]; // @[rawFloatFromFN.scala 47:23]
  wire [9:0] mulAddRecFN_io_b_rawIn_fractIn = io_b[9:0]; // @[rawFloatFromFN.scala 48:25]
  wire  mulAddRecFN_io_b_rawIn_isZeroExpIn = mulAddRecFN_io_b_rawIn_expIn == 5'h0; // @[rawFloatFromFN.scala 50:34]
  wire  mulAddRecFN_io_b_rawIn_isZeroFractIn = mulAddRecFN_io_b_rawIn_fractIn == 10'h0; // @[rawFloatFromFN.scala 51:38]
  wire [3:0] _mulAddRecFN_io_b_rawIn_normDist_T_10 = mulAddRecFN_io_b_rawIn_fractIn[1] ? 4'h8 : 4'h9; // @[Mux.scala 47:69]
  wire [3:0] _mulAddRecFN_io_b_rawIn_normDist_T_11 = mulAddRecFN_io_b_rawIn_fractIn[2] ? 4'h7 :
    _mulAddRecFN_io_b_rawIn_normDist_T_10; // @[Mux.scala 47:69]
  wire [3:0] _mulAddRecFN_io_b_rawIn_normDist_T_12 = mulAddRecFN_io_b_rawIn_fractIn[3] ? 4'h6 :
    _mulAddRecFN_io_b_rawIn_normDist_T_11; // @[Mux.scala 47:69]
  wire [3:0] _mulAddRecFN_io_b_rawIn_normDist_T_13 = mulAddRecFN_io_b_rawIn_fractIn[4] ? 4'h5 :
    _mulAddRecFN_io_b_rawIn_normDist_T_12; // @[Mux.scala 47:69]
  wire [3:0] _mulAddRecFN_io_b_rawIn_normDist_T_14 = mulAddRecFN_io_b_rawIn_fractIn[5] ? 4'h4 :
    _mulAddRecFN_io_b_rawIn_normDist_T_13; // @[Mux.scala 47:69]
  wire [3:0] _mulAddRecFN_io_b_rawIn_normDist_T_15 = mulAddRecFN_io_b_rawIn_fractIn[6] ? 4'h3 :
    _mulAddRecFN_io_b_rawIn_normDist_T_14; // @[Mux.scala 47:69]
  wire [3:0] _mulAddRecFN_io_b_rawIn_normDist_T_16 = mulAddRecFN_io_b_rawIn_fractIn[7] ? 4'h2 :
    _mulAddRecFN_io_b_rawIn_normDist_T_15; // @[Mux.scala 47:69]
  wire [3:0] _mulAddRecFN_io_b_rawIn_normDist_T_17 = mulAddRecFN_io_b_rawIn_fractIn[8] ? 4'h1 :
    _mulAddRecFN_io_b_rawIn_normDist_T_16; // @[Mux.scala 47:69]
  wire [3:0] mulAddRecFN_io_b_rawIn_normDist = mulAddRecFN_io_b_rawIn_fractIn[9] ? 4'h0 :
    _mulAddRecFN_io_b_rawIn_normDist_T_17; // @[Mux.scala 47:69]
  wire [24:0] _GEN_5 = {{15'd0}, mulAddRecFN_io_b_rawIn_fractIn}; // @[rawFloatFromFN.scala 54:36]
  wire [24:0] _mulAddRecFN_io_b_rawIn_subnormFract_T = _GEN_5 << mulAddRecFN_io_b_rawIn_normDist; // @[rawFloatFromFN.scala 54:36]
  wire [9:0] mulAddRecFN_io_b_rawIn_subnormFract = {_mulAddRecFN_io_b_rawIn_subnormFract_T[8:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  wire [5:0] _GEN_6 = {{2'd0}, mulAddRecFN_io_b_rawIn_normDist}; // @[rawFloatFromFN.scala 57:26]
  wire [5:0] _mulAddRecFN_io_b_rawIn_adjustedExp_T = _GEN_6 ^ 6'h3f; // @[rawFloatFromFN.scala 57:26]
  wire [5:0] _mulAddRecFN_io_b_rawIn_adjustedExp_T_1 = mulAddRecFN_io_b_rawIn_isZeroExpIn ?
    _mulAddRecFN_io_b_rawIn_adjustedExp_T : {{1'd0}, mulAddRecFN_io_b_rawIn_expIn}; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _mulAddRecFN_io_b_rawIn_adjustedExp_T_2 = mulAddRecFN_io_b_rawIn_isZeroExpIn ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  wire [4:0] _GEN_7 = {{3'd0}, _mulAddRecFN_io_b_rawIn_adjustedExp_T_2}; // @[rawFloatFromFN.scala 60:22]
  wire [4:0] _mulAddRecFN_io_b_rawIn_adjustedExp_T_3 = 5'h10 | _GEN_7; // @[rawFloatFromFN.scala 60:22]
  wire [5:0] _GEN_8 = {{1'd0}, _mulAddRecFN_io_b_rawIn_adjustedExp_T_3}; // @[rawFloatFromFN.scala 59:15]
  wire [5:0] mulAddRecFN_io_b_rawIn_adjustedExp = _mulAddRecFN_io_b_rawIn_adjustedExp_T_1 + _GEN_8; // @[rawFloatFromFN.scala 59:15]
  wire  mulAddRecFN_io_b_rawIn_isZero = mulAddRecFN_io_b_rawIn_isZeroExpIn & mulAddRecFN_io_b_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 62:34]
  wire  mulAddRecFN_io_b_rawIn_isSpecial = mulAddRecFN_io_b_rawIn_adjustedExp[5:4] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  wire  mulAddRecFN_io_b_rawIn__isNaN = mulAddRecFN_io_b_rawIn_isSpecial & ~mulAddRecFN_io_b_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 66:33]
  wire [6:0] mulAddRecFN_io_b_rawIn__sExp = {1'b0,$signed(mulAddRecFN_io_b_rawIn_adjustedExp)}; // @[rawFloatFromFN.scala 70:48]
  wire  mulAddRecFN_io_b_rawIn_out_sig_hi_lo = ~mulAddRecFN_io_b_rawIn_isZero; // @[rawFloatFromFN.scala 72:29]
  wire [9:0] mulAddRecFN_io_b_rawIn_out_sig_lo = mulAddRecFN_io_b_rawIn_isZeroExpIn ?
    mulAddRecFN_io_b_rawIn_subnormFract : mulAddRecFN_io_b_rawIn_fractIn; // @[rawFloatFromFN.scala 72:42]
  wire [11:0] mulAddRecFN_io_b_rawIn__sig = {1'h0,mulAddRecFN_io_b_rawIn_out_sig_hi_lo,mulAddRecFN_io_b_rawIn_out_sig_lo
    }; // @[Cat.scala 30:58]
  wire [2:0] _mulAddRecFN_io_b_T_1 = mulAddRecFN_io_b_rawIn_isZero ? 3'h0 : mulAddRecFN_io_b_rawIn__sExp[5:3]; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_9 = {{2'd0}, mulAddRecFN_io_b_rawIn__isNaN}; // @[recFNFromFN.scala 48:79]
  wire [2:0] mulAddRecFN_io_b_hi_lo = _mulAddRecFN_io_b_T_1 | _GEN_9; // @[recFNFromFN.scala 48:79]
  wire [2:0] mulAddRecFN_io_b_lo_hi = mulAddRecFN_io_b_rawIn__sExp[2:0]; // @[recFNFromFN.scala 50:23]
  wire [9:0] mulAddRecFN_io_b_lo_lo = mulAddRecFN_io_b_rawIn__sig[9:0]; // @[recFNFromFN.scala 51:22]
  wire [12:0] mulAddRecFN_io_b_lo = {mulAddRecFN_io_b_lo_hi,mulAddRecFN_io_b_lo_lo}; // @[Cat.scala 30:58]
  wire [3:0] mulAddRecFN_io_b_hi = {mulAddRecFN_io_b_rawIn_sign,mulAddRecFN_io_b_hi_lo}; // @[Cat.scala 30:58]
  wire  mulAddRecFN_io_c_rawIn_sign = io_c[15]; // @[rawFloatFromFN.scala 46:22]
  wire [4:0] mulAddRecFN_io_c_rawIn_expIn = io_c[14:10]; // @[rawFloatFromFN.scala 47:23]
  wire [9:0] mulAddRecFN_io_c_rawIn_fractIn = io_c[9:0]; // @[rawFloatFromFN.scala 48:25]
  wire  mulAddRecFN_io_c_rawIn_isZeroExpIn = mulAddRecFN_io_c_rawIn_expIn == 5'h0; // @[rawFloatFromFN.scala 50:34]
  wire  mulAddRecFN_io_c_rawIn_isZeroFractIn = mulAddRecFN_io_c_rawIn_fractIn == 10'h0; // @[rawFloatFromFN.scala 51:38]
  wire [3:0] _mulAddRecFN_io_c_rawIn_normDist_T_10 = mulAddRecFN_io_c_rawIn_fractIn[1] ? 4'h8 : 4'h9; // @[Mux.scala 47:69]
  wire [3:0] _mulAddRecFN_io_c_rawIn_normDist_T_11 = mulAddRecFN_io_c_rawIn_fractIn[2] ? 4'h7 :
    _mulAddRecFN_io_c_rawIn_normDist_T_10; // @[Mux.scala 47:69]
  wire [3:0] _mulAddRecFN_io_c_rawIn_normDist_T_12 = mulAddRecFN_io_c_rawIn_fractIn[3] ? 4'h6 :
    _mulAddRecFN_io_c_rawIn_normDist_T_11; // @[Mux.scala 47:69]
  wire [3:0] _mulAddRecFN_io_c_rawIn_normDist_T_13 = mulAddRecFN_io_c_rawIn_fractIn[4] ? 4'h5 :
    _mulAddRecFN_io_c_rawIn_normDist_T_12; // @[Mux.scala 47:69]
  wire [3:0] _mulAddRecFN_io_c_rawIn_normDist_T_14 = mulAddRecFN_io_c_rawIn_fractIn[5] ? 4'h4 :
    _mulAddRecFN_io_c_rawIn_normDist_T_13; // @[Mux.scala 47:69]
  wire [3:0] _mulAddRecFN_io_c_rawIn_normDist_T_15 = mulAddRecFN_io_c_rawIn_fractIn[6] ? 4'h3 :
    _mulAddRecFN_io_c_rawIn_normDist_T_14; // @[Mux.scala 47:69]
  wire [3:0] _mulAddRecFN_io_c_rawIn_normDist_T_16 = mulAddRecFN_io_c_rawIn_fractIn[7] ? 4'h2 :
    _mulAddRecFN_io_c_rawIn_normDist_T_15; // @[Mux.scala 47:69]
  wire [3:0] _mulAddRecFN_io_c_rawIn_normDist_T_17 = mulAddRecFN_io_c_rawIn_fractIn[8] ? 4'h1 :
    _mulAddRecFN_io_c_rawIn_normDist_T_16; // @[Mux.scala 47:69]
  wire [3:0] mulAddRecFN_io_c_rawIn_normDist = mulAddRecFN_io_c_rawIn_fractIn[9] ? 4'h0 :
    _mulAddRecFN_io_c_rawIn_normDist_T_17; // @[Mux.scala 47:69]
  wire [24:0] _GEN_10 = {{15'd0}, mulAddRecFN_io_c_rawIn_fractIn}; // @[rawFloatFromFN.scala 54:36]
  wire [24:0] _mulAddRecFN_io_c_rawIn_subnormFract_T = _GEN_10 << mulAddRecFN_io_c_rawIn_normDist; // @[rawFloatFromFN.scala 54:36]
  wire [9:0] mulAddRecFN_io_c_rawIn_subnormFract = {_mulAddRecFN_io_c_rawIn_subnormFract_T[8:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  wire [5:0] _GEN_11 = {{2'd0}, mulAddRecFN_io_c_rawIn_normDist}; // @[rawFloatFromFN.scala 57:26]
  wire [5:0] _mulAddRecFN_io_c_rawIn_adjustedExp_T = _GEN_11 ^ 6'h3f; // @[rawFloatFromFN.scala 57:26]
  wire [5:0] _mulAddRecFN_io_c_rawIn_adjustedExp_T_1 = mulAddRecFN_io_c_rawIn_isZeroExpIn ?
    _mulAddRecFN_io_c_rawIn_adjustedExp_T : {{1'd0}, mulAddRecFN_io_c_rawIn_expIn}; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _mulAddRecFN_io_c_rawIn_adjustedExp_T_2 = mulAddRecFN_io_c_rawIn_isZeroExpIn ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  wire [4:0] _GEN_12 = {{3'd0}, _mulAddRecFN_io_c_rawIn_adjustedExp_T_2}; // @[rawFloatFromFN.scala 60:22]
  wire [4:0] _mulAddRecFN_io_c_rawIn_adjustedExp_T_3 = 5'h10 | _GEN_12; // @[rawFloatFromFN.scala 60:22]
  wire [5:0] _GEN_13 = {{1'd0}, _mulAddRecFN_io_c_rawIn_adjustedExp_T_3}; // @[rawFloatFromFN.scala 59:15]
  wire [5:0] mulAddRecFN_io_c_rawIn_adjustedExp = _mulAddRecFN_io_c_rawIn_adjustedExp_T_1 + _GEN_13; // @[rawFloatFromFN.scala 59:15]
  wire  mulAddRecFN_io_c_rawIn_isZero = mulAddRecFN_io_c_rawIn_isZeroExpIn & mulAddRecFN_io_c_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 62:34]
  wire  mulAddRecFN_io_c_rawIn_isSpecial = mulAddRecFN_io_c_rawIn_adjustedExp[5:4] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  wire  mulAddRecFN_io_c_rawIn__isNaN = mulAddRecFN_io_c_rawIn_isSpecial & ~mulAddRecFN_io_c_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 66:33]
  wire [6:0] mulAddRecFN_io_c_rawIn__sExp = {1'b0,$signed(mulAddRecFN_io_c_rawIn_adjustedExp)}; // @[rawFloatFromFN.scala 70:48]
  wire  mulAddRecFN_io_c_rawIn_out_sig_hi_lo = ~mulAddRecFN_io_c_rawIn_isZero; // @[rawFloatFromFN.scala 72:29]
  wire [9:0] mulAddRecFN_io_c_rawIn_out_sig_lo = mulAddRecFN_io_c_rawIn_isZeroExpIn ?
    mulAddRecFN_io_c_rawIn_subnormFract : mulAddRecFN_io_c_rawIn_fractIn; // @[rawFloatFromFN.scala 72:42]
  wire [11:0] mulAddRecFN_io_c_rawIn__sig = {1'h0,mulAddRecFN_io_c_rawIn_out_sig_hi_lo,mulAddRecFN_io_c_rawIn_out_sig_lo
    }; // @[Cat.scala 30:58]
  wire [2:0] _mulAddRecFN_io_c_T_1 = mulAddRecFN_io_c_rawIn_isZero ? 3'h0 : mulAddRecFN_io_c_rawIn__sExp[5:3]; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_14 = {{2'd0}, mulAddRecFN_io_c_rawIn__isNaN}; // @[recFNFromFN.scala 48:79]
  wire [2:0] mulAddRecFN_io_c_hi_lo = _mulAddRecFN_io_c_T_1 | _GEN_14; // @[recFNFromFN.scala 48:79]
  wire [2:0] mulAddRecFN_io_c_lo_hi = mulAddRecFN_io_c_rawIn__sExp[2:0]; // @[recFNFromFN.scala 50:23]
  wire [9:0] mulAddRecFN_io_c_lo_lo = mulAddRecFN_io_c_rawIn__sig[9:0]; // @[recFNFromFN.scala 51:22]
  wire [12:0] mulAddRecFN_io_c_lo = {mulAddRecFN_io_c_lo_hi,mulAddRecFN_io_c_lo_lo}; // @[Cat.scala 30:58]
  wire [3:0] mulAddRecFN_io_c_hi = {mulAddRecFN_io_c_rawIn_sign,mulAddRecFN_io_c_hi_lo}; // @[Cat.scala 30:58]
  wire [5:0] io_out_rawIn_exp = mulAddRecFN_io_out[15:10]; // @[rawFloatFromRecFN.scala 50:21]
  wire  io_out_rawIn_isZero = io_out_rawIn_exp[5:3] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  wire  io_out_rawIn_isSpecial = io_out_rawIn_exp[5:4] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  wire  io_out_rawIn__isNaN = io_out_rawIn_isSpecial & io_out_rawIn_exp[3]; // @[rawFloatFromRecFN.scala 55:33]
  wire  io_out_rawIn__isInf = io_out_rawIn_isSpecial & ~io_out_rawIn_exp[3]; // @[rawFloatFromRecFN.scala 56:33]
  wire  io_out_rawIn__sign = mulAddRecFN_io_out[16]; // @[rawFloatFromRecFN.scala 58:25]
  wire [6:0] io_out_rawIn__sExp = {1'b0,$signed(io_out_rawIn_exp)}; // @[rawFloatFromRecFN.scala 59:27]
  wire  io_out_rawIn_out_sig_hi_lo = ~io_out_rawIn_isZero; // @[rawFloatFromRecFN.scala 60:39]
  wire [9:0] io_out_rawIn_out_sig_lo = mulAddRecFN_io_out[9:0]; // @[rawFloatFromRecFN.scala 60:51]
  wire [11:0] io_out_rawIn__sig = {1'h0,io_out_rawIn_out_sig_hi_lo,io_out_rawIn_out_sig_lo}; // @[Cat.scala 30:58]
  wire  io_out_isSubnormal = $signed(io_out_rawIn__sExp) < 7'sh12; // @[fNFromRecFN.scala 51:39]
  wire [3:0] io_out_denormShiftDist = 4'h1 - io_out_rawIn__sExp[3:0]; // @[fNFromRecFN.scala 52:39]
  wire [10:0] _io_out_denormFract_T_1 = io_out_rawIn__sig[11:1] >> io_out_denormShiftDist; // @[fNFromRecFN.scala 53:42]
  wire [9:0] io_out_denormFract = _io_out_denormFract_T_1[9:0]; // @[fNFromRecFN.scala 53:60]
  wire [4:0] _io_out_expOut_T_2 = io_out_rawIn__sExp[4:0] - 5'h11; // @[fNFromRecFN.scala 58:45]
  wire [4:0] _io_out_expOut_T_3 = io_out_isSubnormal ? 5'h0 : _io_out_expOut_T_2; // @[fNFromRecFN.scala 56:16]
  wire  _io_out_expOut_T_4 = io_out_rawIn__isNaN | io_out_rawIn__isInf; // @[fNFromRecFN.scala 60:44]
  wire [4:0] _io_out_expOut_T_6 = _io_out_expOut_T_4 ? 5'h1f : 5'h0; // @[Bitwise.scala 72:12]
  wire [4:0] io_out_hi_lo = _io_out_expOut_T_3 | _io_out_expOut_T_6; // @[fNFromRecFN.scala 60:15]
  wire [9:0] _io_out_fractOut_T_1 = io_out_rawIn__isInf ? 10'h0 : io_out_rawIn__sig[9:0]; // @[fNFromRecFN.scala 64:20]
  wire [9:0] io_out_lo = io_out_isSubnormal ? io_out_denormFract : _io_out_fractOut_T_1; // @[fNFromRecFN.scala 62:16]
  wire [5:0] io_out_hi = {io_out_rawIn__sign,io_out_hi_lo}; // @[Cat.scala 30:58]
  MulAddRecFN mulAddRecFN ( // @[hardfloat.scala 31:29]
    .io_a(mulAddRecFN_io_a),
    .io_b(mulAddRecFN_io_b),
    .io_c(mulAddRecFN_io_c),
    .io_out(mulAddRecFN_io_out),
    .io_mulOut(mulAddRecFN_io_mulOut),
    .io_mulIn1(mulAddRecFN_io_mulIn1),
    .io_mulIn2(mulAddRecFN_io_mulIn2),
    .io_correctMulOut(mulAddRecFN_io_correctMulOut),
    .io_correctMulIn(mulAddRecFN_io_correctMulIn),
    .io_sigSum_Msb(mulAddRecFN_io_sigSum_Msb)
  );
  assign io_out = {io_out_hi,io_out_lo}; // @[Cat.scala 30:58]
  assign mulAddRecFN_io_a = {mulAddRecFN_io_a_hi,mulAddRecFN_io_a_lo}; // @[Cat.scala 30:58]
  assign mulAddRecFN_io_b = {mulAddRecFN_io_b_hi,mulAddRecFN_io_b_lo}; // @[Cat.scala 30:58]
  assign mulAddRecFN_io_c = {mulAddRecFN_io_c_hi,mulAddRecFN_io_c_lo}; // @[Cat.scala 30:58]
endmodule
module PE(
  input         clock,
  input         reset,
  input  [15:0] io_FromAbovePE,
  input  [15:0] io_FromL1,
  input  [11:0] io_control_signal_mask,
  output [15:0] io_ToRightPE,
  output [15:0] io_ToBelowPE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] FP16MAC_io_a; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_b; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_c; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_out; // @[PEArray.scala 72:23]
  reg [5:0] L0Index; // @[PEArray.scala 39:24]
  reg [15:0] L0Memory_0; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_1; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_2; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_3; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_4; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_5; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_6; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_7; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_8; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_9; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_10; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_11; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_12; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_13; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_14; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_15; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_16; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_17; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_18; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_19; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_20; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_21; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_22; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_23; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_24; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_25; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_26; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_27; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_28; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_29; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_30; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_31; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_32; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_33; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_34; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_35; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_36; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_37; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_38; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_39; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_40; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_41; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_42; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_43; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_44; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_45; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_46; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_47; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_48; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_49; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_50; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_51; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_52; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_53; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_54; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_55; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_56; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_57; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_58; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_59; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_60; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_61; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_62; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_63; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_64; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_65; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_66; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_67; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_68; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_69; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_70; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_71; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_72; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_73; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_74; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_75; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_76; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_77; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_78; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_79; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_80; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_81; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_82; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_83; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_84; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_85; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_86; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_87; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_88; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_89; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_90; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_91; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_92; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_93; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_94; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_95; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_96; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_97; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_98; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_99; // @[PEArray.scala 40:21]
  reg [2:0] state; // @[PEArray.scala 100:22]
  wire  _T_3 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_12 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_16 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_22 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_31 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_41 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_342 = _T_41 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 231:12 PEArray.scala 32:8]
  wire  _GEN_349 = _T_31 ? 1'h0 : _GEN_342; // @[Conditional.scala 39:67 PEArray.scala 208:12]
  wire  _GEN_459 = _T_22 | _GEN_349; // @[Conditional.scala 39:67 PEArray.scala 32:8]
  wire  _GEN_463 = _T_16 ? 1'h0 : _GEN_459; // @[Conditional.scala 39:67]
  wire  _GEN_572 = _T_12 | _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 149:12]
  wire  sel1 = _T_3 | _GEN_572; // @[Conditional.scala 40:58 PEArray.scala 108:12]
  wire [15:0] MAC_out = FP16MAC_io_out; // @[PEArray.scala 47:21 PEArray.scala 85:11]
  wire  _GEN_465 = _T_16 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 177:12]
  wire  _GEN_580 = _T_12 | _GEN_465; // @[Conditional.scala 39:67 PEArray.scala 34:8]
  wire  sel3 = _T_3 | _GEN_580; // @[Conditional.scala 40:58 PEArray.scala 110:12]
  wire [1:0] _GEN_344 = _T_41 ? 2'h2 : 2'h0; // @[Conditional.scala 39:67 PEArray.scala 233:12 PEArray.scala 35:8]
  wire [1:0] _GEN_351 = _T_31 ? 2'h2 : _GEN_344; // @[Conditional.scala 39:67 PEArray.scala 210:12]
  wire [1:0] _GEN_461 = _T_22 ? 2'h0 : _GEN_351; // @[Conditional.scala 39:67 PEArray.scala 35:8]
  wire [1:0] _GEN_466 = _T_16 ? 2'h0 : _GEN_461; // @[Conditional.scala 39:67 PEArray.scala 178:12]
  wire [1:0] _GEN_574 = _T_12 ? 2'h0 : _GEN_466; // @[Conditional.scala 39:67]
  wire [1:0] sel4 = _T_3 ? 2'h0 : _GEN_574; // @[Conditional.scala 40:58 PEArray.scala 111:12]
  wire [15:0] _GEN_3 = sel4 == 2'h2 ? io_FromL1 : 16'h0; // @[PEArray.scala 65:28 PEArray.scala 66:15 PEArray.scala 69:15]
  wire [15:0] _GEN_4 = sel4 == 2'h1 ? io_FromAbovePE : _GEN_3; // @[PEArray.scala 62:28 PEArray.scala 63:15]
  wire [15:0] mux4out = sel4 == 2'h0 ? 16'h0 : _GEN_4; // @[PEArray.scala 59:22 PEArray.scala 60:13]
  wire [15:0] _GEN_7 = 6'h1 == L0Index ? L0Memory_1 : L0Memory_0; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_8 = 6'h2 == L0Index ? L0Memory_2 : _GEN_7; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_9 = 6'h3 == L0Index ? L0Memory_3 : _GEN_8; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_10 = 6'h4 == L0Index ? L0Memory_4 : _GEN_9; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_11 = 6'h5 == L0Index ? L0Memory_5 : _GEN_10; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_12 = 6'h6 == L0Index ? L0Memory_6 : _GEN_11; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_13 = 6'h7 == L0Index ? L0Memory_7 : _GEN_12; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_14 = 6'h8 == L0Index ? L0Memory_8 : _GEN_13; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_15 = 6'h9 == L0Index ? L0Memory_9 : _GEN_14; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_16 = 6'ha == L0Index ? L0Memory_10 : _GEN_15; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_17 = 6'hb == L0Index ? L0Memory_11 : _GEN_16; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_18 = 6'hc == L0Index ? L0Memory_12 : _GEN_17; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_19 = 6'hd == L0Index ? L0Memory_13 : _GEN_18; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_20 = 6'he == L0Index ? L0Memory_14 : _GEN_19; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_21 = 6'hf == L0Index ? L0Memory_15 : _GEN_20; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_22 = 6'h10 == L0Index ? L0Memory_16 : _GEN_21; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_23 = 6'h11 == L0Index ? L0Memory_17 : _GEN_22; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_24 = 6'h12 == L0Index ? L0Memory_18 : _GEN_23; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_25 = 6'h13 == L0Index ? L0Memory_19 : _GEN_24; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_26 = 6'h14 == L0Index ? L0Memory_20 : _GEN_25; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_27 = 6'h15 == L0Index ? L0Memory_21 : _GEN_26; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_28 = 6'h16 == L0Index ? L0Memory_22 : _GEN_27; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_29 = 6'h17 == L0Index ? L0Memory_23 : _GEN_28; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_30 = 6'h18 == L0Index ? L0Memory_24 : _GEN_29; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_31 = 6'h19 == L0Index ? L0Memory_25 : _GEN_30; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_32 = 6'h1a == L0Index ? L0Memory_26 : _GEN_31; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_33 = 6'h1b == L0Index ? L0Memory_27 : _GEN_32; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_34 = 6'h1c == L0Index ? L0Memory_28 : _GEN_33; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_35 = 6'h1d == L0Index ? L0Memory_29 : _GEN_34; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_36 = 6'h1e == L0Index ? L0Memory_30 : _GEN_35; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_37 = 6'h1f == L0Index ? L0Memory_31 : _GEN_36; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_38 = 6'h20 == L0Index ? L0Memory_32 : _GEN_37; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_39 = 6'h21 == L0Index ? L0Memory_33 : _GEN_38; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_40 = 6'h22 == L0Index ? L0Memory_34 : _GEN_39; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_41 = 6'h23 == L0Index ? L0Memory_35 : _GEN_40; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_42 = 6'h24 == L0Index ? L0Memory_36 : _GEN_41; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_43 = 6'h25 == L0Index ? L0Memory_37 : _GEN_42; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_44 = 6'h26 == L0Index ? L0Memory_38 : _GEN_43; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_45 = 6'h27 == L0Index ? L0Memory_39 : _GEN_44; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_46 = 6'h28 == L0Index ? L0Memory_40 : _GEN_45; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_47 = 6'h29 == L0Index ? L0Memory_41 : _GEN_46; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_48 = 6'h2a == L0Index ? L0Memory_42 : _GEN_47; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_49 = 6'h2b == L0Index ? L0Memory_43 : _GEN_48; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_50 = 6'h2c == L0Index ? L0Memory_44 : _GEN_49; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_51 = 6'h2d == L0Index ? L0Memory_45 : _GEN_50; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_52 = 6'h2e == L0Index ? L0Memory_46 : _GEN_51; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_53 = 6'h2f == L0Index ? L0Memory_47 : _GEN_52; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_54 = 6'h30 == L0Index ? L0Memory_48 : _GEN_53; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_55 = 6'h31 == L0Index ? L0Memory_49 : _GEN_54; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_56 = 6'h32 == L0Index ? L0Memory_50 : _GEN_55; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_57 = 6'h33 == L0Index ? L0Memory_51 : _GEN_56; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_58 = 6'h34 == L0Index ? L0Memory_52 : _GEN_57; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_59 = 6'h35 == L0Index ? L0Memory_53 : _GEN_58; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_60 = 6'h36 == L0Index ? L0Memory_54 : _GEN_59; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_61 = 6'h37 == L0Index ? L0Memory_55 : _GEN_60; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_62 = 6'h38 == L0Index ? L0Memory_56 : _GEN_61; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_63 = 6'h39 == L0Index ? L0Memory_57 : _GEN_62; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_64 = 6'h3a == L0Index ? L0Memory_58 : _GEN_63; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_65 = 6'h3b == L0Index ? L0Memory_59 : _GEN_64; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_66 = 6'h3c == L0Index ? L0Memory_60 : _GEN_65; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_67 = 6'h3d == L0Index ? L0Memory_61 : _GEN_66; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_68 = 6'h3e == L0Index ? L0Memory_62 : _GEN_67; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_69 = 6'h3f == L0Index ? L0Memory_63 : _GEN_68; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [6:0] _GEN_793 = {{1'd0}, L0Index}; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_70 = 7'h40 == _GEN_793 ? L0Memory_64 : _GEN_69; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_71 = 7'h41 == _GEN_793 ? L0Memory_65 : _GEN_70; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_72 = 7'h42 == _GEN_793 ? L0Memory_66 : _GEN_71; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_73 = 7'h43 == _GEN_793 ? L0Memory_67 : _GEN_72; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_74 = 7'h44 == _GEN_793 ? L0Memory_68 : _GEN_73; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_75 = 7'h45 == _GEN_793 ? L0Memory_69 : _GEN_74; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_76 = 7'h46 == _GEN_793 ? L0Memory_70 : _GEN_75; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_77 = 7'h47 == _GEN_793 ? L0Memory_71 : _GEN_76; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_78 = 7'h48 == _GEN_793 ? L0Memory_72 : _GEN_77; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_79 = 7'h49 == _GEN_793 ? L0Memory_73 : _GEN_78; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_80 = 7'h4a == _GEN_793 ? L0Memory_74 : _GEN_79; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_81 = 7'h4b == _GEN_793 ? L0Memory_75 : _GEN_80; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_82 = 7'h4c == _GEN_793 ? L0Memory_76 : _GEN_81; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_83 = 7'h4d == _GEN_793 ? L0Memory_77 : _GEN_82; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_84 = 7'h4e == _GEN_793 ? L0Memory_78 : _GEN_83; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_85 = 7'h4f == _GEN_793 ? L0Memory_79 : _GEN_84; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_86 = 7'h50 == _GEN_793 ? L0Memory_80 : _GEN_85; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_87 = 7'h51 == _GEN_793 ? L0Memory_81 : _GEN_86; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_88 = 7'h52 == _GEN_793 ? L0Memory_82 : _GEN_87; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_89 = 7'h53 == _GEN_793 ? L0Memory_83 : _GEN_88; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_90 = 7'h54 == _GEN_793 ? L0Memory_84 : _GEN_89; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_91 = 7'h55 == _GEN_793 ? L0Memory_85 : _GEN_90; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_92 = 7'h56 == _GEN_793 ? L0Memory_86 : _GEN_91; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_93 = 7'h57 == _GEN_793 ? L0Memory_87 : _GEN_92; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_94 = 7'h58 == _GEN_793 ? L0Memory_88 : _GEN_93; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_95 = 7'h59 == _GEN_793 ? L0Memory_89 : _GEN_94; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_96 = 7'h5a == _GEN_793 ? L0Memory_90 : _GEN_95; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_97 = 7'h5b == _GEN_793 ? L0Memory_91 : _GEN_96; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_98 = 7'h5c == _GEN_793 ? L0Memory_92 : _GEN_97; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_99 = 7'h5d == _GEN_793 ? L0Memory_93 : _GEN_98; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_100 = 7'h5e == _GEN_793 ? L0Memory_94 : _GEN_99; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_101 = 7'h5f == _GEN_793 ? L0Memory_95 : _GEN_100; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_102 = 7'h60 == _GEN_793 ? L0Memory_96 : _GEN_101; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_103 = 7'h61 == _GEN_793 ? L0Memory_97 : _GEN_102; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_104 = 7'h62 == _GEN_793 ? L0Memory_98 : _GEN_103; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_105 = 7'h63 == _GEN_793 ? L0Memory_99 : _GEN_104; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire  _GEN_575 = _T_12 ? 1'h0 : _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 157:12]
  wire  sel5 = _T_3 ? 1'h0 : _GEN_575; // @[Conditional.scala 40:58 PEArray.scala 112:12]
  reg [15:0] mux2out_reg; // @[PEArray.scala 90:28]
  reg [15:0] mux3out_reg; // @[PEArray.scala 91:28]
  reg [9:0] count; // @[PEArray.scala 101:22]
  reg [5:0] GRU_out_width; // @[PEArray.scala 104:26]
  wire [7:0] _GEN_118 = io_control_signal_mask[11] ? 8'h0 : {{2'd0}, GRU_out_width}; // @[PEArray.scala 116:57 PEArray.scala 145:23 PEArray.scala 104:26]
  wire [9:0] _count_T_1 = count + 10'h1; // @[PEArray.scala 162:24]
  wire [9:0] _GEN_120 = count != 10'h33 ? _count_T_1 : count; // @[PEArray.scala 161:27 PEArray.scala 162:15 PEArray.scala 101:22]
  wire [9:0] _GEN_124 = count != 10'h188 ? _count_T_1 : count; // @[PEArray.scala 183:28 PEArray.scala 184:15 PEArray.scala 101:22]
  wire [9:0] _GEN_125 = count == 10'h188 ? 10'h0 : _GEN_124; // @[PEArray.scala 186:28 PEArray.scala 187:15]
  wire [2:0] _GEN_126 = count == 10'h188 ? 3'h0 : state; // @[PEArray.scala 186:28 PEArray.scala 188:15 PEArray.scala 100:22]
  wire [9:0] _GEN_127 = count != 10'h0 ? _count_T_1 : count; // @[PEArray.scala 192:32 PEArray.scala 193:15 PEArray.scala 101:22]
  wire  _T_24 = count == 10'h0; // @[PEArray.scala 195:18]
  wire [5:0] _GEN_128 = count == 10'h0 ? 6'h0 : L0Index; // @[PEArray.scala 195:26 PEArray.scala 196:17 PEArray.scala 39:24]
  wire [9:0] _T_27 = 10'h0 - 10'h1; // @[PEArray.scala 198:51]
  wire [15:0] _GEN_129 = 6'h0 == L0Index ? io_FromL1 : L0Memory_0; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_130 = 6'h1 == L0Index ? io_FromL1 : L0Memory_1; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_131 = 6'h2 == L0Index ? io_FromL1 : L0Memory_2; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_132 = 6'h3 == L0Index ? io_FromL1 : L0Memory_3; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_133 = 6'h4 == L0Index ? io_FromL1 : L0Memory_4; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_134 = 6'h5 == L0Index ? io_FromL1 : L0Memory_5; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_135 = 6'h6 == L0Index ? io_FromL1 : L0Memory_6; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_136 = 6'h7 == L0Index ? io_FromL1 : L0Memory_7; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_137 = 6'h8 == L0Index ? io_FromL1 : L0Memory_8; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_138 = 6'h9 == L0Index ? io_FromL1 : L0Memory_9; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_139 = 6'ha == L0Index ? io_FromL1 : L0Memory_10; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_140 = 6'hb == L0Index ? io_FromL1 : L0Memory_11; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_141 = 6'hc == L0Index ? io_FromL1 : L0Memory_12; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_142 = 6'hd == L0Index ? io_FromL1 : L0Memory_13; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_143 = 6'he == L0Index ? io_FromL1 : L0Memory_14; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_144 = 6'hf == L0Index ? io_FromL1 : L0Memory_15; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_145 = 6'h10 == L0Index ? io_FromL1 : L0Memory_16; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_146 = 6'h11 == L0Index ? io_FromL1 : L0Memory_17; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_147 = 6'h12 == L0Index ? io_FromL1 : L0Memory_18; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_148 = 6'h13 == L0Index ? io_FromL1 : L0Memory_19; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_149 = 6'h14 == L0Index ? io_FromL1 : L0Memory_20; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_150 = 6'h15 == L0Index ? io_FromL1 : L0Memory_21; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_151 = 6'h16 == L0Index ? io_FromL1 : L0Memory_22; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_152 = 6'h17 == L0Index ? io_FromL1 : L0Memory_23; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_153 = 6'h18 == L0Index ? io_FromL1 : L0Memory_24; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_154 = 6'h19 == L0Index ? io_FromL1 : L0Memory_25; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_155 = 6'h1a == L0Index ? io_FromL1 : L0Memory_26; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_156 = 6'h1b == L0Index ? io_FromL1 : L0Memory_27; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_157 = 6'h1c == L0Index ? io_FromL1 : L0Memory_28; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_158 = 6'h1d == L0Index ? io_FromL1 : L0Memory_29; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_159 = 6'h1e == L0Index ? io_FromL1 : L0Memory_30; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_160 = 6'h1f == L0Index ? io_FromL1 : L0Memory_31; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_161 = 6'h20 == L0Index ? io_FromL1 : L0Memory_32; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_162 = 6'h21 == L0Index ? io_FromL1 : L0Memory_33; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_163 = 6'h22 == L0Index ? io_FromL1 : L0Memory_34; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_164 = 6'h23 == L0Index ? io_FromL1 : L0Memory_35; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_165 = 6'h24 == L0Index ? io_FromL1 : L0Memory_36; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_166 = 6'h25 == L0Index ? io_FromL1 : L0Memory_37; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_167 = 6'h26 == L0Index ? io_FromL1 : L0Memory_38; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_168 = 6'h27 == L0Index ? io_FromL1 : L0Memory_39; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_169 = 6'h28 == L0Index ? io_FromL1 : L0Memory_40; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_170 = 6'h29 == L0Index ? io_FromL1 : L0Memory_41; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_171 = 6'h2a == L0Index ? io_FromL1 : L0Memory_42; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_172 = 6'h2b == L0Index ? io_FromL1 : L0Memory_43; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_173 = 6'h2c == L0Index ? io_FromL1 : L0Memory_44; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_174 = 6'h2d == L0Index ? io_FromL1 : L0Memory_45; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_175 = 6'h2e == L0Index ? io_FromL1 : L0Memory_46; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_176 = 6'h2f == L0Index ? io_FromL1 : L0Memory_47; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_177 = 6'h30 == L0Index ? io_FromL1 : L0Memory_48; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_178 = 6'h31 == L0Index ? io_FromL1 : L0Memory_49; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_179 = 6'h32 == L0Index ? io_FromL1 : L0Memory_50; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_180 = 6'h33 == L0Index ? io_FromL1 : L0Memory_51; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_181 = 6'h34 == L0Index ? io_FromL1 : L0Memory_52; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_182 = 6'h35 == L0Index ? io_FromL1 : L0Memory_53; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_183 = 6'h36 == L0Index ? io_FromL1 : L0Memory_54; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_184 = 6'h37 == L0Index ? io_FromL1 : L0Memory_55; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_185 = 6'h38 == L0Index ? io_FromL1 : L0Memory_56; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_186 = 6'h39 == L0Index ? io_FromL1 : L0Memory_57; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_187 = 6'h3a == L0Index ? io_FromL1 : L0Memory_58; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_188 = 6'h3b == L0Index ? io_FromL1 : L0Memory_59; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_189 = 6'h3c == L0Index ? io_FromL1 : L0Memory_60; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_190 = 6'h3d == L0Index ? io_FromL1 : L0Memory_61; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_191 = 6'h3e == L0Index ? io_FromL1 : L0Memory_62; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_192 = 6'h3f == L0Index ? io_FromL1 : L0Memory_63; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_193 = 7'h40 == _GEN_793 ? io_FromL1 : L0Memory_64; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_194 = 7'h41 == _GEN_793 ? io_FromL1 : L0Memory_65; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_195 = 7'h42 == _GEN_793 ? io_FromL1 : L0Memory_66; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_196 = 7'h43 == _GEN_793 ? io_FromL1 : L0Memory_67; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_197 = 7'h44 == _GEN_793 ? io_FromL1 : L0Memory_68; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_198 = 7'h45 == _GEN_793 ? io_FromL1 : L0Memory_69; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_199 = 7'h46 == _GEN_793 ? io_FromL1 : L0Memory_70; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_200 = 7'h47 == _GEN_793 ? io_FromL1 : L0Memory_71; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_201 = 7'h48 == _GEN_793 ? io_FromL1 : L0Memory_72; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_202 = 7'h49 == _GEN_793 ? io_FromL1 : L0Memory_73; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_203 = 7'h4a == _GEN_793 ? io_FromL1 : L0Memory_74; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_204 = 7'h4b == _GEN_793 ? io_FromL1 : L0Memory_75; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_205 = 7'h4c == _GEN_793 ? io_FromL1 : L0Memory_76; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_206 = 7'h4d == _GEN_793 ? io_FromL1 : L0Memory_77; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_207 = 7'h4e == _GEN_793 ? io_FromL1 : L0Memory_78; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_208 = 7'h4f == _GEN_793 ? io_FromL1 : L0Memory_79; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_209 = 7'h50 == _GEN_793 ? io_FromL1 : L0Memory_80; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_210 = 7'h51 == _GEN_793 ? io_FromL1 : L0Memory_81; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_211 = 7'h52 == _GEN_793 ? io_FromL1 : L0Memory_82; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_212 = 7'h53 == _GEN_793 ? io_FromL1 : L0Memory_83; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_213 = 7'h54 == _GEN_793 ? io_FromL1 : L0Memory_84; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_214 = 7'h55 == _GEN_793 ? io_FromL1 : L0Memory_85; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_215 = 7'h56 == _GEN_793 ? io_FromL1 : L0Memory_86; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_216 = 7'h57 == _GEN_793 ? io_FromL1 : L0Memory_87; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_217 = 7'h58 == _GEN_793 ? io_FromL1 : L0Memory_88; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_218 = 7'h59 == _GEN_793 ? io_FromL1 : L0Memory_89; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_219 = 7'h5a == _GEN_793 ? io_FromL1 : L0Memory_90; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_220 = 7'h5b == _GEN_793 ? io_FromL1 : L0Memory_91; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_221 = 7'h5c == _GEN_793 ? io_FromL1 : L0Memory_92; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_222 = 7'h5d == _GEN_793 ? io_FromL1 : L0Memory_93; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_223 = 7'h5e == _GEN_793 ? io_FromL1 : L0Memory_94; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_224 = 7'h5f == _GEN_793 ? io_FromL1 : L0Memory_95; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_225 = 7'h60 == _GEN_793 ? io_FromL1 : L0Memory_96; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_226 = 7'h61 == _GEN_793 ? io_FromL1 : L0Memory_97; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_227 = 7'h62 == _GEN_793 ? io_FromL1 : L0Memory_98; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_228 = 7'h63 == _GEN_793 ? io_FromL1 : L0Memory_99; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [5:0] _L0Index_T_2 = L0Index + 6'h1; // @[PEArray.scala 200:28]
  wire [15:0] _GEN_229 = count >= 10'h1 & count <= _T_27 ? _GEN_129 : L0Memory_0; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_230 = count >= 10'h1 & count <= _T_27 ? _GEN_130 : L0Memory_1; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_231 = count >= 10'h1 & count <= _T_27 ? _GEN_131 : L0Memory_2; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_232 = count >= 10'h1 & count <= _T_27 ? _GEN_132 : L0Memory_3; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_233 = count >= 10'h1 & count <= _T_27 ? _GEN_133 : L0Memory_4; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_234 = count >= 10'h1 & count <= _T_27 ? _GEN_134 : L0Memory_5; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_235 = count >= 10'h1 & count <= _T_27 ? _GEN_135 : L0Memory_6; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_236 = count >= 10'h1 & count <= _T_27 ? _GEN_136 : L0Memory_7; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_237 = count >= 10'h1 & count <= _T_27 ? _GEN_137 : L0Memory_8; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_238 = count >= 10'h1 & count <= _T_27 ? _GEN_138 : L0Memory_9; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_239 = count >= 10'h1 & count <= _T_27 ? _GEN_139 : L0Memory_10; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_240 = count >= 10'h1 & count <= _T_27 ? _GEN_140 : L0Memory_11; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_241 = count >= 10'h1 & count <= _T_27 ? _GEN_141 : L0Memory_12; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_242 = count >= 10'h1 & count <= _T_27 ? _GEN_142 : L0Memory_13; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_243 = count >= 10'h1 & count <= _T_27 ? _GEN_143 : L0Memory_14; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_244 = count >= 10'h1 & count <= _T_27 ? _GEN_144 : L0Memory_15; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_245 = count >= 10'h1 & count <= _T_27 ? _GEN_145 : L0Memory_16; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_246 = count >= 10'h1 & count <= _T_27 ? _GEN_146 : L0Memory_17; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_247 = count >= 10'h1 & count <= _T_27 ? _GEN_147 : L0Memory_18; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_248 = count >= 10'h1 & count <= _T_27 ? _GEN_148 : L0Memory_19; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_249 = count >= 10'h1 & count <= _T_27 ? _GEN_149 : L0Memory_20; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_250 = count >= 10'h1 & count <= _T_27 ? _GEN_150 : L0Memory_21; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_251 = count >= 10'h1 & count <= _T_27 ? _GEN_151 : L0Memory_22; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_252 = count >= 10'h1 & count <= _T_27 ? _GEN_152 : L0Memory_23; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_253 = count >= 10'h1 & count <= _T_27 ? _GEN_153 : L0Memory_24; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_254 = count >= 10'h1 & count <= _T_27 ? _GEN_154 : L0Memory_25; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_255 = count >= 10'h1 & count <= _T_27 ? _GEN_155 : L0Memory_26; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_256 = count >= 10'h1 & count <= _T_27 ? _GEN_156 : L0Memory_27; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_257 = count >= 10'h1 & count <= _T_27 ? _GEN_157 : L0Memory_28; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_258 = count >= 10'h1 & count <= _T_27 ? _GEN_158 : L0Memory_29; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_259 = count >= 10'h1 & count <= _T_27 ? _GEN_159 : L0Memory_30; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_260 = count >= 10'h1 & count <= _T_27 ? _GEN_160 : L0Memory_31; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_261 = count >= 10'h1 & count <= _T_27 ? _GEN_161 : L0Memory_32; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_262 = count >= 10'h1 & count <= _T_27 ? _GEN_162 : L0Memory_33; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_263 = count >= 10'h1 & count <= _T_27 ? _GEN_163 : L0Memory_34; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_264 = count >= 10'h1 & count <= _T_27 ? _GEN_164 : L0Memory_35; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_265 = count >= 10'h1 & count <= _T_27 ? _GEN_165 : L0Memory_36; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_266 = count >= 10'h1 & count <= _T_27 ? _GEN_166 : L0Memory_37; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_267 = count >= 10'h1 & count <= _T_27 ? _GEN_167 : L0Memory_38; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_268 = count >= 10'h1 & count <= _T_27 ? _GEN_168 : L0Memory_39; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_269 = count >= 10'h1 & count <= _T_27 ? _GEN_169 : L0Memory_40; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_270 = count >= 10'h1 & count <= _T_27 ? _GEN_170 : L0Memory_41; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_271 = count >= 10'h1 & count <= _T_27 ? _GEN_171 : L0Memory_42; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_272 = count >= 10'h1 & count <= _T_27 ? _GEN_172 : L0Memory_43; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_273 = count >= 10'h1 & count <= _T_27 ? _GEN_173 : L0Memory_44; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_274 = count >= 10'h1 & count <= _T_27 ? _GEN_174 : L0Memory_45; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_275 = count >= 10'h1 & count <= _T_27 ? _GEN_175 : L0Memory_46; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_276 = count >= 10'h1 & count <= _T_27 ? _GEN_176 : L0Memory_47; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_277 = count >= 10'h1 & count <= _T_27 ? _GEN_177 : L0Memory_48; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_278 = count >= 10'h1 & count <= _T_27 ? _GEN_178 : L0Memory_49; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_279 = count >= 10'h1 & count <= _T_27 ? _GEN_179 : L0Memory_50; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_280 = count >= 10'h1 & count <= _T_27 ? _GEN_180 : L0Memory_51; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_281 = count >= 10'h1 & count <= _T_27 ? _GEN_181 : L0Memory_52; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_282 = count >= 10'h1 & count <= _T_27 ? _GEN_182 : L0Memory_53; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_283 = count >= 10'h1 & count <= _T_27 ? _GEN_183 : L0Memory_54; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_284 = count >= 10'h1 & count <= _T_27 ? _GEN_184 : L0Memory_55; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_285 = count >= 10'h1 & count <= _T_27 ? _GEN_185 : L0Memory_56; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_286 = count >= 10'h1 & count <= _T_27 ? _GEN_186 : L0Memory_57; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_287 = count >= 10'h1 & count <= _T_27 ? _GEN_187 : L0Memory_58; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_288 = count >= 10'h1 & count <= _T_27 ? _GEN_188 : L0Memory_59; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_289 = count >= 10'h1 & count <= _T_27 ? _GEN_189 : L0Memory_60; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_290 = count >= 10'h1 & count <= _T_27 ? _GEN_190 : L0Memory_61; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_291 = count >= 10'h1 & count <= _T_27 ? _GEN_191 : L0Memory_62; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_292 = count >= 10'h1 & count <= _T_27 ? _GEN_192 : L0Memory_63; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_293 = count >= 10'h1 & count <= _T_27 ? _GEN_193 : L0Memory_64; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_294 = count >= 10'h1 & count <= _T_27 ? _GEN_194 : L0Memory_65; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_295 = count >= 10'h1 & count <= _T_27 ? _GEN_195 : L0Memory_66; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_296 = count >= 10'h1 & count <= _T_27 ? _GEN_196 : L0Memory_67; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_297 = count >= 10'h1 & count <= _T_27 ? _GEN_197 : L0Memory_68; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_298 = count >= 10'h1 & count <= _T_27 ? _GEN_198 : L0Memory_69; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_299 = count >= 10'h1 & count <= _T_27 ? _GEN_199 : L0Memory_70; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_300 = count >= 10'h1 & count <= _T_27 ? _GEN_200 : L0Memory_71; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_301 = count >= 10'h1 & count <= _T_27 ? _GEN_201 : L0Memory_72; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_302 = count >= 10'h1 & count <= _T_27 ? _GEN_202 : L0Memory_73; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_303 = count >= 10'h1 & count <= _T_27 ? _GEN_203 : L0Memory_74; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_304 = count >= 10'h1 & count <= _T_27 ? _GEN_204 : L0Memory_75; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_305 = count >= 10'h1 & count <= _T_27 ? _GEN_205 : L0Memory_76; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_306 = count >= 10'h1 & count <= _T_27 ? _GEN_206 : L0Memory_77; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_307 = count >= 10'h1 & count <= _T_27 ? _GEN_207 : L0Memory_78; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_308 = count >= 10'h1 & count <= _T_27 ? _GEN_208 : L0Memory_79; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_309 = count >= 10'h1 & count <= _T_27 ? _GEN_209 : L0Memory_80; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_310 = count >= 10'h1 & count <= _T_27 ? _GEN_210 : L0Memory_81; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_311 = count >= 10'h1 & count <= _T_27 ? _GEN_211 : L0Memory_82; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_312 = count >= 10'h1 & count <= _T_27 ? _GEN_212 : L0Memory_83; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_313 = count >= 10'h1 & count <= _T_27 ? _GEN_213 : L0Memory_84; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_314 = count >= 10'h1 & count <= _T_27 ? _GEN_214 : L0Memory_85; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_315 = count >= 10'h1 & count <= _T_27 ? _GEN_215 : L0Memory_86; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_316 = count >= 10'h1 & count <= _T_27 ? _GEN_216 : L0Memory_87; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_317 = count >= 10'h1 & count <= _T_27 ? _GEN_217 : L0Memory_88; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_318 = count >= 10'h1 & count <= _T_27 ? _GEN_218 : L0Memory_89; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_319 = count >= 10'h1 & count <= _T_27 ? _GEN_219 : L0Memory_90; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_320 = count >= 10'h1 & count <= _T_27 ? _GEN_220 : L0Memory_91; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_321 = count >= 10'h1 & count <= _T_27 ? _GEN_221 : L0Memory_92; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_322 = count >= 10'h1 & count <= _T_27 ? _GEN_222 : L0Memory_93; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_323 = count >= 10'h1 & count <= _T_27 ? _GEN_223 : L0Memory_94; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_324 = count >= 10'h1 & count <= _T_27 ? _GEN_224 : L0Memory_95; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_325 = count >= 10'h1 & count <= _T_27 ? _GEN_225 : L0Memory_96; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_326 = count >= 10'h1 & count <= _T_27 ? _GEN_226 : L0Memory_97; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_327 = count >= 10'h1 & count <= _T_27 ? _GEN_227 : L0Memory_98; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_328 = count >= 10'h1 & count <= _T_27 ? _GEN_228 : L0Memory_99; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [5:0] _GEN_329 = count >= 10'h1 & count <= _T_27 ? _L0Index_T_2 : _GEN_128; // @[PEArray.scala 198:59 PEArray.scala 200:17]
  wire [9:0] _GEN_330 = _T_24 ? 10'h0 : _GEN_127; // @[PEArray.scala 202:32 PEArray.scala 203:15]
  wire [2:0] _GEN_331 = _T_24 ? 3'h0 : state; // @[PEArray.scala 202:32 PEArray.scala 204:15 PEArray.scala 100:22]
  wire [9:0] _GEN_865 = {{4'd0}, GRU_out_width}; // @[PEArray.scala 220:19]
  wire [9:0] _GEN_0 = count % _GEN_865; // @[PEArray.scala 220:19]
  wire [5:0] _T_36 = _GEN_0[5:0]; // @[PEArray.scala 220:19]
  wire [5:0] _T_38 = GRU_out_width - 6'h1; // @[PEArray.scala 220:55]
  wire [5:0] _GEN_334 = _T_36 == _T_38 ? _L0Index_T_2 : 6'h0; // @[PEArray.scala 220:62 PEArray.scala 221:17 PEArray.scala 214:15]
  wire [5:0] _GEN_346 = _T_41 ? _GEN_334 : L0Index; // @[Conditional.scala 39:67 PEArray.scala 39:24]
  wire [9:0] _GEN_347 = _T_41 ? _GEN_330 : count; // @[Conditional.scala 39:67 PEArray.scala 101:22]
  wire [2:0] _GEN_348 = _T_41 ? _GEN_331 : state; // @[Conditional.scala 39:67 PEArray.scala 100:22]
  wire [5:0] _GEN_353 = _T_31 ? _GEN_334 : _GEN_346; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_354 = _T_31 ? _GEN_330 : _GEN_347; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_355 = _T_31 ? _GEN_331 : _GEN_348; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_356 = _T_22 ? _GEN_330 : _GEN_354; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_357 = _T_22 ? _GEN_329 : _GEN_353; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_458 = _T_22 ? _GEN_331 : _GEN_355; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_690 = _T_3 ? _GEN_118 : {{2'd0}, GRU_out_width}; // @[Conditional.scala 40:58 PEArray.scala 104:26]
  FP16MulAdder FP16MAC ( // @[PEArray.scala 72:23]
    .io_a(FP16MAC_io_a),
    .io_b(FP16MAC_io_b),
    .io_c(FP16MAC_io_c),
    .io_out(FP16MAC_io_out)
  );
  assign io_ToRightPE = mux3out_reg; // @[PEArray.scala 95:16]
  assign io_ToBelowPE = mux2out_reg; // @[PEArray.scala 94:16]
  assign FP16MAC_io_a = sel1 ? io_FromL1 : 16'h0; // @[PEArray.scala 50:14 PEArray.scala 50:23 PEArray.scala 51:24]
  assign FP16MAC_io_b = sel5 ? mux4out : _GEN_105; // @[PEArray.scala 77:13 PEArray.scala 78:18 PEArray.scala 81:18]
  assign FP16MAC_io_c = sel5 ? _GEN_105 : mux4out; // @[PEArray.scala 77:13 PEArray.scala 79:18 PEArray.scala 82:18]
  always @(posedge clock) begin
    if (reset) begin // @[PEArray.scala 39:24]
      L0Index <= 6'h0; // @[PEArray.scala 39:24]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h0; // @[PEArray.scala 159:15]
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h3; // @[PEArray.scala 181:15]
      end else begin
        L0Index <= _GEN_357;
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_0 <= _GEN_229;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_1 <= _GEN_230;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_2 <= _GEN_231;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_3 <= _GEN_232;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_4 <= _GEN_233;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_5 <= _GEN_234;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_6 <= _GEN_235;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_7 <= _GEN_236;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_8 <= _GEN_237;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_9 <= _GEN_238;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_10 <= _GEN_239;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_11 <= _GEN_240;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_12 <= _GEN_241;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_13 <= _GEN_242;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_14 <= _GEN_243;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_15 <= _GEN_244;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_16 <= _GEN_245;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_17 <= _GEN_246;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_18 <= _GEN_247;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_19 <= _GEN_248;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_20 <= _GEN_249;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_21 <= _GEN_250;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_22 <= _GEN_251;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_23 <= _GEN_252;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_24 <= _GEN_253;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_25 <= _GEN_254;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_26 <= _GEN_255;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_27 <= _GEN_256;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_28 <= _GEN_257;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_29 <= _GEN_258;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_30 <= _GEN_259;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_31 <= _GEN_260;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_32 <= _GEN_261;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_33 <= _GEN_262;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_34 <= _GEN_263;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_35 <= _GEN_264;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_36 <= _GEN_265;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_37 <= _GEN_266;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_38 <= _GEN_267;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_39 <= _GEN_268;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_40 <= _GEN_269;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_41 <= _GEN_270;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_42 <= _GEN_271;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_43 <= _GEN_272;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_44 <= _GEN_273;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_45 <= _GEN_274;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_46 <= _GEN_275;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_47 <= _GEN_276;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_48 <= _GEN_277;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_49 <= _GEN_278;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_50 <= _GEN_279;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_51 <= _GEN_280;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_52 <= _GEN_281;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_53 <= _GEN_282;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_54 <= _GEN_283;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_55 <= _GEN_284;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_56 <= _GEN_285;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_57 <= _GEN_286;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_58 <= _GEN_287;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_59 <= _GEN_288;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_60 <= _GEN_289;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_61 <= _GEN_290;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_62 <= _GEN_291;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_63 <= _GEN_292;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_64 <= _GEN_293;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_65 <= _GEN_294;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_66 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_67 <= _GEN_296;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_68 <= _GEN_297;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_69 <= _GEN_298;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_70 <= _GEN_299;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_71 <= _GEN_300;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_72 <= _GEN_301;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_73 <= _GEN_302;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_74 <= _GEN_303;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_75 <= _GEN_304;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_76 <= _GEN_305;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_77 <= _GEN_306;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_78 <= _GEN_307;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_79 <= _GEN_308;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_80 <= _GEN_309;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_81 <= _GEN_310;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_82 <= _GEN_311;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_83 <= _GEN_312;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_84 <= _GEN_313;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_85 <= _GEN_314;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_86 <= _GEN_315;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_87 <= _GEN_316;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_88 <= _GEN_317;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_89 <= _GEN_318;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_90 <= _GEN_319;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_91 <= _GEN_320;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_92 <= _GEN_321;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_93 <= _GEN_322;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_94 <= _GEN_323;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_95 <= _GEN_324;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_96 <= _GEN_325;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_97 <= _GEN_326;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_98 <= _GEN_327;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_99 <= _GEN_328;
          end
        end
      end
    end
    if (reset) begin // @[PEArray.scala 100:22]
      state <= 3'h0; // @[PEArray.scala 100:22]
    end else if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[11]) begin // @[PEArray.scala 116:57]
        state <= 3'h1;
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      if (count == 10'h33) begin // @[PEArray.scala 164:27]
        state <= 3'h0; // @[PEArray.scala 166:15]
      end
    end else if (_T_16) begin // @[Conditional.scala 39:67]
      state <= _GEN_126;
    end else begin
      state <= _GEN_458;
    end
    if (reset) begin // @[PEArray.scala 90:28]
      mux2out_reg <= 16'h0; // @[PEArray.scala 90:28]
    end else begin
      mux2out_reg <= MAC_out; // @[PEArray.scala 90:28]
    end
    if (reset) begin // @[PEArray.scala 91:28]
      mux3out_reg <= 16'h0; // @[PEArray.scala 91:28]
    end else if (sel3) begin // @[PEArray.scala 56:14]
      mux3out_reg <= MAC_out; // @[PEArray.scala 56:23]
    end else if (sel1) begin // @[PEArray.scala 50:14]
      mux3out_reg <= io_FromL1; // @[PEArray.scala 50:23]
    end else begin
      mux3out_reg <= 16'h0; // @[PEArray.scala 51:24]
    end
    if (reset) begin // @[PEArray.scala 101:22]
      count <= 10'h0; // @[PEArray.scala 101:22]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        if (count == 10'h33) begin // @[PEArray.scala 164:27]
          count <= 10'h0; // @[PEArray.scala 165:15]
        end else begin
          count <= _GEN_120;
        end
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        count <= _GEN_125;
      end else begin
        count <= _GEN_356;
      end
    end
    GRU_out_width <= _GEN_690[5:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  L0Index = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  L0Memory_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  L0Memory_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  L0Memory_2 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  L0Memory_3 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  L0Memory_4 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  L0Memory_5 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  L0Memory_6 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  L0Memory_7 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  L0Memory_8 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  L0Memory_9 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  L0Memory_10 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  L0Memory_11 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  L0Memory_12 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  L0Memory_13 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  L0Memory_14 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  L0Memory_15 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  L0Memory_16 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  L0Memory_17 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  L0Memory_18 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  L0Memory_19 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  L0Memory_20 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  L0Memory_21 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  L0Memory_22 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  L0Memory_23 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  L0Memory_24 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  L0Memory_25 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  L0Memory_26 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  L0Memory_27 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  L0Memory_28 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  L0Memory_29 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  L0Memory_30 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  L0Memory_31 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  L0Memory_32 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  L0Memory_33 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  L0Memory_34 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  L0Memory_35 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  L0Memory_36 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  L0Memory_37 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  L0Memory_38 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  L0Memory_39 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  L0Memory_40 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  L0Memory_41 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  L0Memory_42 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  L0Memory_43 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  L0Memory_44 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  L0Memory_45 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  L0Memory_46 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  L0Memory_47 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  L0Memory_48 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  L0Memory_49 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  L0Memory_50 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  L0Memory_51 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  L0Memory_52 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  L0Memory_53 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  L0Memory_54 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  L0Memory_55 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  L0Memory_56 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  L0Memory_57 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  L0Memory_58 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  L0Memory_59 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  L0Memory_60 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  L0Memory_61 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  L0Memory_62 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  L0Memory_63 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  L0Memory_64 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  L0Memory_65 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  L0Memory_66 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  L0Memory_67 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  L0Memory_68 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  L0Memory_69 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  L0Memory_70 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  L0Memory_71 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  L0Memory_72 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  L0Memory_73 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  L0Memory_74 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  L0Memory_75 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  L0Memory_76 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  L0Memory_77 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  L0Memory_78 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  L0Memory_79 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  L0Memory_80 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  L0Memory_81 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  L0Memory_82 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  L0Memory_83 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  L0Memory_84 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  L0Memory_85 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  L0Memory_86 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  L0Memory_87 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  L0Memory_88 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  L0Memory_89 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  L0Memory_90 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  L0Memory_91 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  L0Memory_92 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  L0Memory_93 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  L0Memory_94 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  L0Memory_95 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  L0Memory_96 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  L0Memory_97 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  L0Memory_98 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  L0Memory_99 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  state = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  mux2out_reg = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  mux3out_reg = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  count = _RAND_104[9:0];
  _RAND_105 = {1{`RANDOM}};
  GRU_out_width = _RAND_105[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PE_1(
  input         clock,
  input         reset,
  input  [15:0] io_FromAbovePE,
  input  [15:0] io_FromL1,
  input  [11:0] io_control_signal_mask,
  output [15:0] io_ToRightPE,
  output [15:0] io_ToBelowPE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] FP16MAC_io_a; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_b; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_c; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_out; // @[PEArray.scala 72:23]
  reg [5:0] L0Index; // @[PEArray.scala 39:24]
  reg [15:0] L0Memory_0; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_1; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_2; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_3; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_4; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_5; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_6; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_7; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_8; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_9; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_10; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_11; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_12; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_13; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_14; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_15; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_16; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_17; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_18; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_19; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_20; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_21; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_22; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_23; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_24; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_25; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_26; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_27; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_28; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_29; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_30; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_31; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_32; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_33; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_34; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_35; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_36; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_37; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_38; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_39; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_40; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_41; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_42; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_43; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_44; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_45; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_46; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_47; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_48; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_49; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_50; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_51; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_52; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_53; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_54; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_55; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_56; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_57; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_58; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_59; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_60; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_61; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_62; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_63; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_64; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_65; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_66; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_67; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_68; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_69; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_70; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_71; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_72; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_73; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_74; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_75; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_76; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_77; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_78; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_79; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_80; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_81; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_82; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_83; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_84; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_85; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_86; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_87; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_88; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_89; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_90; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_91; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_92; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_93; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_94; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_95; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_96; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_97; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_98; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_99; // @[PEArray.scala 40:21]
  reg [2:0] state; // @[PEArray.scala 100:22]
  wire  _T_3 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_12 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_16 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_22 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_31 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_41 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_342 = _T_41 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 231:12 PEArray.scala 32:8]
  wire  _GEN_349 = _T_31 ? 1'h0 : _GEN_342; // @[Conditional.scala 39:67 PEArray.scala 208:12]
  wire  _GEN_459 = _T_22 | _GEN_349; // @[Conditional.scala 39:67 PEArray.scala 32:8]
  wire  _GEN_463 = _T_16 ? 1'h0 : _GEN_459; // @[Conditional.scala 39:67]
  wire  _GEN_572 = _T_12 | _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 149:12]
  wire  sel1 = _T_3 | _GEN_572; // @[Conditional.scala 40:58 PEArray.scala 108:12]
  wire [15:0] MAC_out = FP16MAC_io_out; // @[PEArray.scala 47:21 PEArray.scala 85:11]
  wire  _GEN_465 = _T_16 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 177:12]
  wire  _GEN_580 = _T_12 | _GEN_465; // @[Conditional.scala 39:67 PEArray.scala 34:8]
  wire  sel3 = _T_3 | _GEN_580; // @[Conditional.scala 40:58 PEArray.scala 110:12]
  wire [1:0] _GEN_344 = _T_41 ? 2'h2 : 2'h0; // @[Conditional.scala 39:67 PEArray.scala 233:12 PEArray.scala 35:8]
  wire [1:0] _GEN_351 = _T_31 ? 2'h2 : _GEN_344; // @[Conditional.scala 39:67 PEArray.scala 210:12]
  wire [1:0] _GEN_461 = _T_22 ? 2'h0 : _GEN_351; // @[Conditional.scala 39:67 PEArray.scala 35:8]
  wire [1:0] _GEN_466 = _T_16 ? 2'h0 : _GEN_461; // @[Conditional.scala 39:67 PEArray.scala 178:12]
  wire [1:0] _GEN_574 = _T_12 ? 2'h1 : _GEN_466; // @[Conditional.scala 39:67]
  wire [1:0] sel4 = _T_3 ? 2'h0 : _GEN_574; // @[Conditional.scala 40:58 PEArray.scala 111:12]
  wire [15:0] _GEN_3 = sel4 == 2'h2 ? io_FromL1 : 16'h0; // @[PEArray.scala 65:28 PEArray.scala 66:15 PEArray.scala 69:15]
  wire [15:0] _GEN_4 = sel4 == 2'h1 ? io_FromAbovePE : _GEN_3; // @[PEArray.scala 62:28 PEArray.scala 63:15]
  wire [15:0] mux4out = sel4 == 2'h0 ? 16'h0 : _GEN_4; // @[PEArray.scala 59:22 PEArray.scala 60:13]
  wire [15:0] _GEN_7 = 6'h1 == L0Index ? L0Memory_1 : L0Memory_0; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_8 = 6'h2 == L0Index ? L0Memory_2 : _GEN_7; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_9 = 6'h3 == L0Index ? L0Memory_3 : _GEN_8; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_10 = 6'h4 == L0Index ? L0Memory_4 : _GEN_9; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_11 = 6'h5 == L0Index ? L0Memory_5 : _GEN_10; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_12 = 6'h6 == L0Index ? L0Memory_6 : _GEN_11; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_13 = 6'h7 == L0Index ? L0Memory_7 : _GEN_12; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_14 = 6'h8 == L0Index ? L0Memory_8 : _GEN_13; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_15 = 6'h9 == L0Index ? L0Memory_9 : _GEN_14; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_16 = 6'ha == L0Index ? L0Memory_10 : _GEN_15; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_17 = 6'hb == L0Index ? L0Memory_11 : _GEN_16; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_18 = 6'hc == L0Index ? L0Memory_12 : _GEN_17; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_19 = 6'hd == L0Index ? L0Memory_13 : _GEN_18; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_20 = 6'he == L0Index ? L0Memory_14 : _GEN_19; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_21 = 6'hf == L0Index ? L0Memory_15 : _GEN_20; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_22 = 6'h10 == L0Index ? L0Memory_16 : _GEN_21; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_23 = 6'h11 == L0Index ? L0Memory_17 : _GEN_22; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_24 = 6'h12 == L0Index ? L0Memory_18 : _GEN_23; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_25 = 6'h13 == L0Index ? L0Memory_19 : _GEN_24; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_26 = 6'h14 == L0Index ? L0Memory_20 : _GEN_25; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_27 = 6'h15 == L0Index ? L0Memory_21 : _GEN_26; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_28 = 6'h16 == L0Index ? L0Memory_22 : _GEN_27; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_29 = 6'h17 == L0Index ? L0Memory_23 : _GEN_28; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_30 = 6'h18 == L0Index ? L0Memory_24 : _GEN_29; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_31 = 6'h19 == L0Index ? L0Memory_25 : _GEN_30; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_32 = 6'h1a == L0Index ? L0Memory_26 : _GEN_31; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_33 = 6'h1b == L0Index ? L0Memory_27 : _GEN_32; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_34 = 6'h1c == L0Index ? L0Memory_28 : _GEN_33; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_35 = 6'h1d == L0Index ? L0Memory_29 : _GEN_34; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_36 = 6'h1e == L0Index ? L0Memory_30 : _GEN_35; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_37 = 6'h1f == L0Index ? L0Memory_31 : _GEN_36; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_38 = 6'h20 == L0Index ? L0Memory_32 : _GEN_37; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_39 = 6'h21 == L0Index ? L0Memory_33 : _GEN_38; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_40 = 6'h22 == L0Index ? L0Memory_34 : _GEN_39; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_41 = 6'h23 == L0Index ? L0Memory_35 : _GEN_40; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_42 = 6'h24 == L0Index ? L0Memory_36 : _GEN_41; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_43 = 6'h25 == L0Index ? L0Memory_37 : _GEN_42; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_44 = 6'h26 == L0Index ? L0Memory_38 : _GEN_43; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_45 = 6'h27 == L0Index ? L0Memory_39 : _GEN_44; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_46 = 6'h28 == L0Index ? L0Memory_40 : _GEN_45; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_47 = 6'h29 == L0Index ? L0Memory_41 : _GEN_46; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_48 = 6'h2a == L0Index ? L0Memory_42 : _GEN_47; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_49 = 6'h2b == L0Index ? L0Memory_43 : _GEN_48; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_50 = 6'h2c == L0Index ? L0Memory_44 : _GEN_49; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_51 = 6'h2d == L0Index ? L0Memory_45 : _GEN_50; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_52 = 6'h2e == L0Index ? L0Memory_46 : _GEN_51; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_53 = 6'h2f == L0Index ? L0Memory_47 : _GEN_52; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_54 = 6'h30 == L0Index ? L0Memory_48 : _GEN_53; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_55 = 6'h31 == L0Index ? L0Memory_49 : _GEN_54; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_56 = 6'h32 == L0Index ? L0Memory_50 : _GEN_55; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_57 = 6'h33 == L0Index ? L0Memory_51 : _GEN_56; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_58 = 6'h34 == L0Index ? L0Memory_52 : _GEN_57; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_59 = 6'h35 == L0Index ? L0Memory_53 : _GEN_58; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_60 = 6'h36 == L0Index ? L0Memory_54 : _GEN_59; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_61 = 6'h37 == L0Index ? L0Memory_55 : _GEN_60; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_62 = 6'h38 == L0Index ? L0Memory_56 : _GEN_61; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_63 = 6'h39 == L0Index ? L0Memory_57 : _GEN_62; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_64 = 6'h3a == L0Index ? L0Memory_58 : _GEN_63; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_65 = 6'h3b == L0Index ? L0Memory_59 : _GEN_64; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_66 = 6'h3c == L0Index ? L0Memory_60 : _GEN_65; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_67 = 6'h3d == L0Index ? L0Memory_61 : _GEN_66; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_68 = 6'h3e == L0Index ? L0Memory_62 : _GEN_67; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_69 = 6'h3f == L0Index ? L0Memory_63 : _GEN_68; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [6:0] _GEN_793 = {{1'd0}, L0Index}; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_70 = 7'h40 == _GEN_793 ? L0Memory_64 : _GEN_69; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_71 = 7'h41 == _GEN_793 ? L0Memory_65 : _GEN_70; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_72 = 7'h42 == _GEN_793 ? L0Memory_66 : _GEN_71; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_73 = 7'h43 == _GEN_793 ? L0Memory_67 : _GEN_72; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_74 = 7'h44 == _GEN_793 ? L0Memory_68 : _GEN_73; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_75 = 7'h45 == _GEN_793 ? L0Memory_69 : _GEN_74; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_76 = 7'h46 == _GEN_793 ? L0Memory_70 : _GEN_75; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_77 = 7'h47 == _GEN_793 ? L0Memory_71 : _GEN_76; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_78 = 7'h48 == _GEN_793 ? L0Memory_72 : _GEN_77; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_79 = 7'h49 == _GEN_793 ? L0Memory_73 : _GEN_78; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_80 = 7'h4a == _GEN_793 ? L0Memory_74 : _GEN_79; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_81 = 7'h4b == _GEN_793 ? L0Memory_75 : _GEN_80; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_82 = 7'h4c == _GEN_793 ? L0Memory_76 : _GEN_81; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_83 = 7'h4d == _GEN_793 ? L0Memory_77 : _GEN_82; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_84 = 7'h4e == _GEN_793 ? L0Memory_78 : _GEN_83; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_85 = 7'h4f == _GEN_793 ? L0Memory_79 : _GEN_84; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_86 = 7'h50 == _GEN_793 ? L0Memory_80 : _GEN_85; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_87 = 7'h51 == _GEN_793 ? L0Memory_81 : _GEN_86; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_88 = 7'h52 == _GEN_793 ? L0Memory_82 : _GEN_87; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_89 = 7'h53 == _GEN_793 ? L0Memory_83 : _GEN_88; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_90 = 7'h54 == _GEN_793 ? L0Memory_84 : _GEN_89; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_91 = 7'h55 == _GEN_793 ? L0Memory_85 : _GEN_90; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_92 = 7'h56 == _GEN_793 ? L0Memory_86 : _GEN_91; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_93 = 7'h57 == _GEN_793 ? L0Memory_87 : _GEN_92; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_94 = 7'h58 == _GEN_793 ? L0Memory_88 : _GEN_93; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_95 = 7'h59 == _GEN_793 ? L0Memory_89 : _GEN_94; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_96 = 7'h5a == _GEN_793 ? L0Memory_90 : _GEN_95; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_97 = 7'h5b == _GEN_793 ? L0Memory_91 : _GEN_96; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_98 = 7'h5c == _GEN_793 ? L0Memory_92 : _GEN_97; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_99 = 7'h5d == _GEN_793 ? L0Memory_93 : _GEN_98; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_100 = 7'h5e == _GEN_793 ? L0Memory_94 : _GEN_99; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_101 = 7'h5f == _GEN_793 ? L0Memory_95 : _GEN_100; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_102 = 7'h60 == _GEN_793 ? L0Memory_96 : _GEN_101; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_103 = 7'h61 == _GEN_793 ? L0Memory_97 : _GEN_102; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_104 = 7'h62 == _GEN_793 ? L0Memory_98 : _GEN_103; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_105 = 7'h63 == _GEN_793 ? L0Memory_99 : _GEN_104; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire  _GEN_575 = _T_12 ? 1'h0 : _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 157:12]
  wire  sel5 = _T_3 ? 1'h0 : _GEN_575; // @[Conditional.scala 40:58 PEArray.scala 112:12]
  reg [15:0] mux2out_reg; // @[PEArray.scala 90:28]
  reg [15:0] mux3out_reg; // @[PEArray.scala 91:28]
  reg [9:0] count; // @[PEArray.scala 101:22]
  reg [5:0] GRU_out_width; // @[PEArray.scala 104:26]
  wire [7:0] _GEN_118 = io_control_signal_mask[11] ? 8'h0 : {{2'd0}, GRU_out_width}; // @[PEArray.scala 116:57 PEArray.scala 145:23 PEArray.scala 104:26]
  wire [9:0] _count_T_1 = count + 10'h1; // @[PEArray.scala 162:24]
  wire [9:0] _GEN_120 = count != 10'h33 ? _count_T_1 : count; // @[PEArray.scala 161:27 PEArray.scala 162:15 PEArray.scala 101:22]
  wire [9:0] _GEN_124 = count != 10'h188 ? _count_T_1 : count; // @[PEArray.scala 183:28 PEArray.scala 184:15 PEArray.scala 101:22]
  wire [9:0] _GEN_125 = count == 10'h188 ? 10'h0 : _GEN_124; // @[PEArray.scala 186:28 PEArray.scala 187:15]
  wire [2:0] _GEN_126 = count == 10'h188 ? 3'h0 : state; // @[PEArray.scala 186:28 PEArray.scala 188:15 PEArray.scala 100:22]
  wire [9:0] _GEN_127 = count != 10'h0 ? _count_T_1 : count; // @[PEArray.scala 192:32 PEArray.scala 193:15 PEArray.scala 101:22]
  wire  _T_24 = count == 10'h0; // @[PEArray.scala 195:18]
  wire [5:0] _GEN_128 = count == 10'h0 ? 6'h0 : L0Index; // @[PEArray.scala 195:26 PEArray.scala 196:17 PEArray.scala 39:24]
  wire [9:0] _T_27 = 10'h0 - 10'h1; // @[PEArray.scala 198:51]
  wire [15:0] _GEN_129 = 6'h0 == L0Index ? io_FromL1 : L0Memory_0; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_130 = 6'h1 == L0Index ? io_FromL1 : L0Memory_1; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_131 = 6'h2 == L0Index ? io_FromL1 : L0Memory_2; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_132 = 6'h3 == L0Index ? io_FromL1 : L0Memory_3; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_133 = 6'h4 == L0Index ? io_FromL1 : L0Memory_4; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_134 = 6'h5 == L0Index ? io_FromL1 : L0Memory_5; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_135 = 6'h6 == L0Index ? io_FromL1 : L0Memory_6; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_136 = 6'h7 == L0Index ? io_FromL1 : L0Memory_7; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_137 = 6'h8 == L0Index ? io_FromL1 : L0Memory_8; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_138 = 6'h9 == L0Index ? io_FromL1 : L0Memory_9; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_139 = 6'ha == L0Index ? io_FromL1 : L0Memory_10; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_140 = 6'hb == L0Index ? io_FromL1 : L0Memory_11; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_141 = 6'hc == L0Index ? io_FromL1 : L0Memory_12; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_142 = 6'hd == L0Index ? io_FromL1 : L0Memory_13; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_143 = 6'he == L0Index ? io_FromL1 : L0Memory_14; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_144 = 6'hf == L0Index ? io_FromL1 : L0Memory_15; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_145 = 6'h10 == L0Index ? io_FromL1 : L0Memory_16; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_146 = 6'h11 == L0Index ? io_FromL1 : L0Memory_17; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_147 = 6'h12 == L0Index ? io_FromL1 : L0Memory_18; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_148 = 6'h13 == L0Index ? io_FromL1 : L0Memory_19; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_149 = 6'h14 == L0Index ? io_FromL1 : L0Memory_20; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_150 = 6'h15 == L0Index ? io_FromL1 : L0Memory_21; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_151 = 6'h16 == L0Index ? io_FromL1 : L0Memory_22; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_152 = 6'h17 == L0Index ? io_FromL1 : L0Memory_23; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_153 = 6'h18 == L0Index ? io_FromL1 : L0Memory_24; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_154 = 6'h19 == L0Index ? io_FromL1 : L0Memory_25; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_155 = 6'h1a == L0Index ? io_FromL1 : L0Memory_26; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_156 = 6'h1b == L0Index ? io_FromL1 : L0Memory_27; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_157 = 6'h1c == L0Index ? io_FromL1 : L0Memory_28; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_158 = 6'h1d == L0Index ? io_FromL1 : L0Memory_29; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_159 = 6'h1e == L0Index ? io_FromL1 : L0Memory_30; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_160 = 6'h1f == L0Index ? io_FromL1 : L0Memory_31; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_161 = 6'h20 == L0Index ? io_FromL1 : L0Memory_32; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_162 = 6'h21 == L0Index ? io_FromL1 : L0Memory_33; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_163 = 6'h22 == L0Index ? io_FromL1 : L0Memory_34; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_164 = 6'h23 == L0Index ? io_FromL1 : L0Memory_35; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_165 = 6'h24 == L0Index ? io_FromL1 : L0Memory_36; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_166 = 6'h25 == L0Index ? io_FromL1 : L0Memory_37; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_167 = 6'h26 == L0Index ? io_FromL1 : L0Memory_38; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_168 = 6'h27 == L0Index ? io_FromL1 : L0Memory_39; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_169 = 6'h28 == L0Index ? io_FromL1 : L0Memory_40; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_170 = 6'h29 == L0Index ? io_FromL1 : L0Memory_41; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_171 = 6'h2a == L0Index ? io_FromL1 : L0Memory_42; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_172 = 6'h2b == L0Index ? io_FromL1 : L0Memory_43; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_173 = 6'h2c == L0Index ? io_FromL1 : L0Memory_44; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_174 = 6'h2d == L0Index ? io_FromL1 : L0Memory_45; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_175 = 6'h2e == L0Index ? io_FromL1 : L0Memory_46; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_176 = 6'h2f == L0Index ? io_FromL1 : L0Memory_47; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_177 = 6'h30 == L0Index ? io_FromL1 : L0Memory_48; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_178 = 6'h31 == L0Index ? io_FromL1 : L0Memory_49; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_179 = 6'h32 == L0Index ? io_FromL1 : L0Memory_50; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_180 = 6'h33 == L0Index ? io_FromL1 : L0Memory_51; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_181 = 6'h34 == L0Index ? io_FromL1 : L0Memory_52; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_182 = 6'h35 == L0Index ? io_FromL1 : L0Memory_53; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_183 = 6'h36 == L0Index ? io_FromL1 : L0Memory_54; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_184 = 6'h37 == L0Index ? io_FromL1 : L0Memory_55; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_185 = 6'h38 == L0Index ? io_FromL1 : L0Memory_56; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_186 = 6'h39 == L0Index ? io_FromL1 : L0Memory_57; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_187 = 6'h3a == L0Index ? io_FromL1 : L0Memory_58; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_188 = 6'h3b == L0Index ? io_FromL1 : L0Memory_59; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_189 = 6'h3c == L0Index ? io_FromL1 : L0Memory_60; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_190 = 6'h3d == L0Index ? io_FromL1 : L0Memory_61; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_191 = 6'h3e == L0Index ? io_FromL1 : L0Memory_62; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_192 = 6'h3f == L0Index ? io_FromL1 : L0Memory_63; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_193 = 7'h40 == _GEN_793 ? io_FromL1 : L0Memory_64; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_194 = 7'h41 == _GEN_793 ? io_FromL1 : L0Memory_65; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_195 = 7'h42 == _GEN_793 ? io_FromL1 : L0Memory_66; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_196 = 7'h43 == _GEN_793 ? io_FromL1 : L0Memory_67; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_197 = 7'h44 == _GEN_793 ? io_FromL1 : L0Memory_68; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_198 = 7'h45 == _GEN_793 ? io_FromL1 : L0Memory_69; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_199 = 7'h46 == _GEN_793 ? io_FromL1 : L0Memory_70; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_200 = 7'h47 == _GEN_793 ? io_FromL1 : L0Memory_71; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_201 = 7'h48 == _GEN_793 ? io_FromL1 : L0Memory_72; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_202 = 7'h49 == _GEN_793 ? io_FromL1 : L0Memory_73; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_203 = 7'h4a == _GEN_793 ? io_FromL1 : L0Memory_74; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_204 = 7'h4b == _GEN_793 ? io_FromL1 : L0Memory_75; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_205 = 7'h4c == _GEN_793 ? io_FromL1 : L0Memory_76; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_206 = 7'h4d == _GEN_793 ? io_FromL1 : L0Memory_77; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_207 = 7'h4e == _GEN_793 ? io_FromL1 : L0Memory_78; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_208 = 7'h4f == _GEN_793 ? io_FromL1 : L0Memory_79; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_209 = 7'h50 == _GEN_793 ? io_FromL1 : L0Memory_80; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_210 = 7'h51 == _GEN_793 ? io_FromL1 : L0Memory_81; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_211 = 7'h52 == _GEN_793 ? io_FromL1 : L0Memory_82; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_212 = 7'h53 == _GEN_793 ? io_FromL1 : L0Memory_83; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_213 = 7'h54 == _GEN_793 ? io_FromL1 : L0Memory_84; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_214 = 7'h55 == _GEN_793 ? io_FromL1 : L0Memory_85; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_215 = 7'h56 == _GEN_793 ? io_FromL1 : L0Memory_86; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_216 = 7'h57 == _GEN_793 ? io_FromL1 : L0Memory_87; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_217 = 7'h58 == _GEN_793 ? io_FromL1 : L0Memory_88; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_218 = 7'h59 == _GEN_793 ? io_FromL1 : L0Memory_89; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_219 = 7'h5a == _GEN_793 ? io_FromL1 : L0Memory_90; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_220 = 7'h5b == _GEN_793 ? io_FromL1 : L0Memory_91; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_221 = 7'h5c == _GEN_793 ? io_FromL1 : L0Memory_92; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_222 = 7'h5d == _GEN_793 ? io_FromL1 : L0Memory_93; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_223 = 7'h5e == _GEN_793 ? io_FromL1 : L0Memory_94; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_224 = 7'h5f == _GEN_793 ? io_FromL1 : L0Memory_95; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_225 = 7'h60 == _GEN_793 ? io_FromL1 : L0Memory_96; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_226 = 7'h61 == _GEN_793 ? io_FromL1 : L0Memory_97; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_227 = 7'h62 == _GEN_793 ? io_FromL1 : L0Memory_98; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_228 = 7'h63 == _GEN_793 ? io_FromL1 : L0Memory_99; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [5:0] _L0Index_T_2 = L0Index + 6'h1; // @[PEArray.scala 200:28]
  wire [15:0] _GEN_229 = count >= 10'h1 & count <= _T_27 ? _GEN_129 : L0Memory_0; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_230 = count >= 10'h1 & count <= _T_27 ? _GEN_130 : L0Memory_1; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_231 = count >= 10'h1 & count <= _T_27 ? _GEN_131 : L0Memory_2; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_232 = count >= 10'h1 & count <= _T_27 ? _GEN_132 : L0Memory_3; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_233 = count >= 10'h1 & count <= _T_27 ? _GEN_133 : L0Memory_4; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_234 = count >= 10'h1 & count <= _T_27 ? _GEN_134 : L0Memory_5; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_235 = count >= 10'h1 & count <= _T_27 ? _GEN_135 : L0Memory_6; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_236 = count >= 10'h1 & count <= _T_27 ? _GEN_136 : L0Memory_7; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_237 = count >= 10'h1 & count <= _T_27 ? _GEN_137 : L0Memory_8; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_238 = count >= 10'h1 & count <= _T_27 ? _GEN_138 : L0Memory_9; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_239 = count >= 10'h1 & count <= _T_27 ? _GEN_139 : L0Memory_10; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_240 = count >= 10'h1 & count <= _T_27 ? _GEN_140 : L0Memory_11; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_241 = count >= 10'h1 & count <= _T_27 ? _GEN_141 : L0Memory_12; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_242 = count >= 10'h1 & count <= _T_27 ? _GEN_142 : L0Memory_13; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_243 = count >= 10'h1 & count <= _T_27 ? _GEN_143 : L0Memory_14; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_244 = count >= 10'h1 & count <= _T_27 ? _GEN_144 : L0Memory_15; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_245 = count >= 10'h1 & count <= _T_27 ? _GEN_145 : L0Memory_16; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_246 = count >= 10'h1 & count <= _T_27 ? _GEN_146 : L0Memory_17; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_247 = count >= 10'h1 & count <= _T_27 ? _GEN_147 : L0Memory_18; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_248 = count >= 10'h1 & count <= _T_27 ? _GEN_148 : L0Memory_19; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_249 = count >= 10'h1 & count <= _T_27 ? _GEN_149 : L0Memory_20; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_250 = count >= 10'h1 & count <= _T_27 ? _GEN_150 : L0Memory_21; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_251 = count >= 10'h1 & count <= _T_27 ? _GEN_151 : L0Memory_22; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_252 = count >= 10'h1 & count <= _T_27 ? _GEN_152 : L0Memory_23; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_253 = count >= 10'h1 & count <= _T_27 ? _GEN_153 : L0Memory_24; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_254 = count >= 10'h1 & count <= _T_27 ? _GEN_154 : L0Memory_25; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_255 = count >= 10'h1 & count <= _T_27 ? _GEN_155 : L0Memory_26; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_256 = count >= 10'h1 & count <= _T_27 ? _GEN_156 : L0Memory_27; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_257 = count >= 10'h1 & count <= _T_27 ? _GEN_157 : L0Memory_28; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_258 = count >= 10'h1 & count <= _T_27 ? _GEN_158 : L0Memory_29; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_259 = count >= 10'h1 & count <= _T_27 ? _GEN_159 : L0Memory_30; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_260 = count >= 10'h1 & count <= _T_27 ? _GEN_160 : L0Memory_31; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_261 = count >= 10'h1 & count <= _T_27 ? _GEN_161 : L0Memory_32; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_262 = count >= 10'h1 & count <= _T_27 ? _GEN_162 : L0Memory_33; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_263 = count >= 10'h1 & count <= _T_27 ? _GEN_163 : L0Memory_34; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_264 = count >= 10'h1 & count <= _T_27 ? _GEN_164 : L0Memory_35; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_265 = count >= 10'h1 & count <= _T_27 ? _GEN_165 : L0Memory_36; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_266 = count >= 10'h1 & count <= _T_27 ? _GEN_166 : L0Memory_37; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_267 = count >= 10'h1 & count <= _T_27 ? _GEN_167 : L0Memory_38; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_268 = count >= 10'h1 & count <= _T_27 ? _GEN_168 : L0Memory_39; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_269 = count >= 10'h1 & count <= _T_27 ? _GEN_169 : L0Memory_40; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_270 = count >= 10'h1 & count <= _T_27 ? _GEN_170 : L0Memory_41; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_271 = count >= 10'h1 & count <= _T_27 ? _GEN_171 : L0Memory_42; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_272 = count >= 10'h1 & count <= _T_27 ? _GEN_172 : L0Memory_43; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_273 = count >= 10'h1 & count <= _T_27 ? _GEN_173 : L0Memory_44; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_274 = count >= 10'h1 & count <= _T_27 ? _GEN_174 : L0Memory_45; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_275 = count >= 10'h1 & count <= _T_27 ? _GEN_175 : L0Memory_46; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_276 = count >= 10'h1 & count <= _T_27 ? _GEN_176 : L0Memory_47; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_277 = count >= 10'h1 & count <= _T_27 ? _GEN_177 : L0Memory_48; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_278 = count >= 10'h1 & count <= _T_27 ? _GEN_178 : L0Memory_49; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_279 = count >= 10'h1 & count <= _T_27 ? _GEN_179 : L0Memory_50; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_280 = count >= 10'h1 & count <= _T_27 ? _GEN_180 : L0Memory_51; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_281 = count >= 10'h1 & count <= _T_27 ? _GEN_181 : L0Memory_52; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_282 = count >= 10'h1 & count <= _T_27 ? _GEN_182 : L0Memory_53; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_283 = count >= 10'h1 & count <= _T_27 ? _GEN_183 : L0Memory_54; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_284 = count >= 10'h1 & count <= _T_27 ? _GEN_184 : L0Memory_55; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_285 = count >= 10'h1 & count <= _T_27 ? _GEN_185 : L0Memory_56; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_286 = count >= 10'h1 & count <= _T_27 ? _GEN_186 : L0Memory_57; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_287 = count >= 10'h1 & count <= _T_27 ? _GEN_187 : L0Memory_58; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_288 = count >= 10'h1 & count <= _T_27 ? _GEN_188 : L0Memory_59; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_289 = count >= 10'h1 & count <= _T_27 ? _GEN_189 : L0Memory_60; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_290 = count >= 10'h1 & count <= _T_27 ? _GEN_190 : L0Memory_61; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_291 = count >= 10'h1 & count <= _T_27 ? _GEN_191 : L0Memory_62; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_292 = count >= 10'h1 & count <= _T_27 ? _GEN_192 : L0Memory_63; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_293 = count >= 10'h1 & count <= _T_27 ? _GEN_193 : L0Memory_64; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_294 = count >= 10'h1 & count <= _T_27 ? _GEN_194 : L0Memory_65; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_295 = count >= 10'h1 & count <= _T_27 ? _GEN_195 : L0Memory_66; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_296 = count >= 10'h1 & count <= _T_27 ? _GEN_196 : L0Memory_67; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_297 = count >= 10'h1 & count <= _T_27 ? _GEN_197 : L0Memory_68; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_298 = count >= 10'h1 & count <= _T_27 ? _GEN_198 : L0Memory_69; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_299 = count >= 10'h1 & count <= _T_27 ? _GEN_199 : L0Memory_70; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_300 = count >= 10'h1 & count <= _T_27 ? _GEN_200 : L0Memory_71; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_301 = count >= 10'h1 & count <= _T_27 ? _GEN_201 : L0Memory_72; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_302 = count >= 10'h1 & count <= _T_27 ? _GEN_202 : L0Memory_73; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_303 = count >= 10'h1 & count <= _T_27 ? _GEN_203 : L0Memory_74; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_304 = count >= 10'h1 & count <= _T_27 ? _GEN_204 : L0Memory_75; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_305 = count >= 10'h1 & count <= _T_27 ? _GEN_205 : L0Memory_76; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_306 = count >= 10'h1 & count <= _T_27 ? _GEN_206 : L0Memory_77; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_307 = count >= 10'h1 & count <= _T_27 ? _GEN_207 : L0Memory_78; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_308 = count >= 10'h1 & count <= _T_27 ? _GEN_208 : L0Memory_79; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_309 = count >= 10'h1 & count <= _T_27 ? _GEN_209 : L0Memory_80; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_310 = count >= 10'h1 & count <= _T_27 ? _GEN_210 : L0Memory_81; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_311 = count >= 10'h1 & count <= _T_27 ? _GEN_211 : L0Memory_82; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_312 = count >= 10'h1 & count <= _T_27 ? _GEN_212 : L0Memory_83; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_313 = count >= 10'h1 & count <= _T_27 ? _GEN_213 : L0Memory_84; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_314 = count >= 10'h1 & count <= _T_27 ? _GEN_214 : L0Memory_85; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_315 = count >= 10'h1 & count <= _T_27 ? _GEN_215 : L0Memory_86; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_316 = count >= 10'h1 & count <= _T_27 ? _GEN_216 : L0Memory_87; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_317 = count >= 10'h1 & count <= _T_27 ? _GEN_217 : L0Memory_88; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_318 = count >= 10'h1 & count <= _T_27 ? _GEN_218 : L0Memory_89; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_319 = count >= 10'h1 & count <= _T_27 ? _GEN_219 : L0Memory_90; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_320 = count >= 10'h1 & count <= _T_27 ? _GEN_220 : L0Memory_91; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_321 = count >= 10'h1 & count <= _T_27 ? _GEN_221 : L0Memory_92; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_322 = count >= 10'h1 & count <= _T_27 ? _GEN_222 : L0Memory_93; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_323 = count >= 10'h1 & count <= _T_27 ? _GEN_223 : L0Memory_94; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_324 = count >= 10'h1 & count <= _T_27 ? _GEN_224 : L0Memory_95; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_325 = count >= 10'h1 & count <= _T_27 ? _GEN_225 : L0Memory_96; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_326 = count >= 10'h1 & count <= _T_27 ? _GEN_226 : L0Memory_97; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_327 = count >= 10'h1 & count <= _T_27 ? _GEN_227 : L0Memory_98; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_328 = count >= 10'h1 & count <= _T_27 ? _GEN_228 : L0Memory_99; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [5:0] _GEN_329 = count >= 10'h1 & count <= _T_27 ? _L0Index_T_2 : _GEN_128; // @[PEArray.scala 198:59 PEArray.scala 200:17]
  wire [9:0] _GEN_330 = _T_24 ? 10'h0 : _GEN_127; // @[PEArray.scala 202:32 PEArray.scala 203:15]
  wire [2:0] _GEN_331 = _T_24 ? 3'h0 : state; // @[PEArray.scala 202:32 PEArray.scala 204:15 PEArray.scala 100:22]
  wire [9:0] _GEN_865 = {{4'd0}, GRU_out_width}; // @[PEArray.scala 220:19]
  wire [9:0] _GEN_0 = count % _GEN_865; // @[PEArray.scala 220:19]
  wire [5:0] _T_36 = _GEN_0[5:0]; // @[PEArray.scala 220:19]
  wire [5:0] _T_38 = GRU_out_width - 6'h1; // @[PEArray.scala 220:55]
  wire [5:0] _GEN_334 = _T_36 == _T_38 ? _L0Index_T_2 : 6'h0; // @[PEArray.scala 220:62 PEArray.scala 221:17 PEArray.scala 214:15]
  wire [5:0] _GEN_346 = _T_41 ? _GEN_334 : L0Index; // @[Conditional.scala 39:67 PEArray.scala 39:24]
  wire [9:0] _GEN_347 = _T_41 ? _GEN_330 : count; // @[Conditional.scala 39:67 PEArray.scala 101:22]
  wire [2:0] _GEN_348 = _T_41 ? _GEN_331 : state; // @[Conditional.scala 39:67 PEArray.scala 100:22]
  wire [5:0] _GEN_353 = _T_31 ? _GEN_334 : _GEN_346; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_354 = _T_31 ? _GEN_330 : _GEN_347; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_355 = _T_31 ? _GEN_331 : _GEN_348; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_356 = _T_22 ? _GEN_330 : _GEN_354; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_357 = _T_22 ? _GEN_329 : _GEN_353; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_458 = _T_22 ? _GEN_331 : _GEN_355; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_690 = _T_3 ? _GEN_118 : {{2'd0}, GRU_out_width}; // @[Conditional.scala 40:58 PEArray.scala 104:26]
  FP16MulAdder FP16MAC ( // @[PEArray.scala 72:23]
    .io_a(FP16MAC_io_a),
    .io_b(FP16MAC_io_b),
    .io_c(FP16MAC_io_c),
    .io_out(FP16MAC_io_out)
  );
  assign io_ToRightPE = mux3out_reg; // @[PEArray.scala 95:16]
  assign io_ToBelowPE = mux2out_reg; // @[PEArray.scala 94:16]
  assign FP16MAC_io_a = sel1 ? io_FromL1 : 16'h0; // @[PEArray.scala 50:14 PEArray.scala 50:23 PEArray.scala 51:24]
  assign FP16MAC_io_b = sel5 ? mux4out : _GEN_105; // @[PEArray.scala 77:13 PEArray.scala 78:18 PEArray.scala 81:18]
  assign FP16MAC_io_c = sel5 ? _GEN_105 : mux4out; // @[PEArray.scala 77:13 PEArray.scala 79:18 PEArray.scala 82:18]
  always @(posedge clock) begin
    if (reset) begin // @[PEArray.scala 39:24]
      L0Index <= 6'h0; // @[PEArray.scala 39:24]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h1; // @[PEArray.scala 159:15]
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h3; // @[PEArray.scala 181:15]
      end else begin
        L0Index <= _GEN_357;
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_0 <= _GEN_229;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_1 <= _GEN_230;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_2 <= _GEN_231;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_3 <= _GEN_232;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_4 <= _GEN_233;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_5 <= _GEN_234;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_6 <= _GEN_235;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_7 <= _GEN_236;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_8 <= _GEN_237;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_9 <= _GEN_238;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_10 <= _GEN_239;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_11 <= _GEN_240;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_12 <= _GEN_241;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_13 <= _GEN_242;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_14 <= _GEN_243;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_15 <= _GEN_244;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_16 <= _GEN_245;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_17 <= _GEN_246;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_18 <= _GEN_247;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_19 <= _GEN_248;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_20 <= _GEN_249;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_21 <= _GEN_250;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_22 <= _GEN_251;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_23 <= _GEN_252;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_24 <= _GEN_253;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_25 <= _GEN_254;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_26 <= _GEN_255;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_27 <= _GEN_256;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_28 <= _GEN_257;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_29 <= _GEN_258;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_30 <= _GEN_259;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_31 <= _GEN_260;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_32 <= _GEN_261;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_33 <= _GEN_262;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_34 <= _GEN_263;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_35 <= _GEN_264;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_36 <= _GEN_265;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_37 <= _GEN_266;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_38 <= _GEN_267;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_39 <= _GEN_268;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_40 <= _GEN_269;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_41 <= _GEN_270;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_42 <= _GEN_271;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_43 <= _GEN_272;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_44 <= _GEN_273;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_45 <= _GEN_274;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_46 <= _GEN_275;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_47 <= _GEN_276;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_48 <= _GEN_277;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_49 <= _GEN_278;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_50 <= _GEN_279;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_51 <= _GEN_280;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_52 <= _GEN_281;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_53 <= _GEN_282;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_54 <= _GEN_283;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_55 <= _GEN_284;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_56 <= _GEN_285;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_57 <= _GEN_286;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_58 <= _GEN_287;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_59 <= _GEN_288;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_60 <= _GEN_289;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_61 <= _GEN_290;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_62 <= _GEN_291;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_63 <= _GEN_292;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_64 <= _GEN_293;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_65 <= _GEN_294;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_66 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_67 <= _GEN_296;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_68 <= _GEN_297;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_69 <= _GEN_298;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_70 <= _GEN_299;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_71 <= _GEN_300;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_72 <= _GEN_301;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_73 <= _GEN_302;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_74 <= _GEN_303;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_75 <= _GEN_304;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_76 <= _GEN_305;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_77 <= _GEN_306;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_78 <= _GEN_307;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_79 <= _GEN_308;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_80 <= _GEN_309;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_81 <= _GEN_310;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_82 <= _GEN_311;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_83 <= _GEN_312;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_84 <= _GEN_313;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_85 <= _GEN_314;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_86 <= _GEN_315;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_87 <= _GEN_316;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_88 <= _GEN_317;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_89 <= _GEN_318;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_90 <= _GEN_319;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_91 <= _GEN_320;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_92 <= _GEN_321;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_93 <= _GEN_322;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_94 <= _GEN_323;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_95 <= _GEN_324;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_96 <= _GEN_325;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_97 <= _GEN_326;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_98 <= _GEN_327;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_99 <= _GEN_328;
          end
        end
      end
    end
    if (reset) begin // @[PEArray.scala 100:22]
      state <= 3'h0; // @[PEArray.scala 100:22]
    end else if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[11]) begin // @[PEArray.scala 116:57]
        state <= 3'h1;
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      if (count == 10'h33) begin // @[PEArray.scala 164:27]
        state <= 3'h0; // @[PEArray.scala 166:15]
      end
    end else if (_T_16) begin // @[Conditional.scala 39:67]
      state <= _GEN_126;
    end else begin
      state <= _GEN_458;
    end
    if (reset) begin // @[PEArray.scala 90:28]
      mux2out_reg <= 16'h0; // @[PEArray.scala 90:28]
    end else begin
      mux2out_reg <= MAC_out; // @[PEArray.scala 90:28]
    end
    if (reset) begin // @[PEArray.scala 91:28]
      mux3out_reg <= 16'h0; // @[PEArray.scala 91:28]
    end else if (sel3) begin // @[PEArray.scala 56:14]
      mux3out_reg <= MAC_out; // @[PEArray.scala 56:23]
    end else if (sel1) begin // @[PEArray.scala 50:14]
      mux3out_reg <= io_FromL1; // @[PEArray.scala 50:23]
    end else begin
      mux3out_reg <= 16'h0; // @[PEArray.scala 51:24]
    end
    if (reset) begin // @[PEArray.scala 101:22]
      count <= 10'h0; // @[PEArray.scala 101:22]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        if (count == 10'h33) begin // @[PEArray.scala 164:27]
          count <= 10'h0; // @[PEArray.scala 165:15]
        end else begin
          count <= _GEN_120;
        end
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        count <= _GEN_125;
      end else begin
        count <= _GEN_356;
      end
    end
    GRU_out_width <= _GEN_690[5:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  L0Index = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  L0Memory_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  L0Memory_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  L0Memory_2 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  L0Memory_3 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  L0Memory_4 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  L0Memory_5 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  L0Memory_6 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  L0Memory_7 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  L0Memory_8 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  L0Memory_9 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  L0Memory_10 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  L0Memory_11 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  L0Memory_12 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  L0Memory_13 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  L0Memory_14 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  L0Memory_15 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  L0Memory_16 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  L0Memory_17 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  L0Memory_18 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  L0Memory_19 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  L0Memory_20 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  L0Memory_21 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  L0Memory_22 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  L0Memory_23 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  L0Memory_24 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  L0Memory_25 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  L0Memory_26 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  L0Memory_27 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  L0Memory_28 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  L0Memory_29 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  L0Memory_30 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  L0Memory_31 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  L0Memory_32 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  L0Memory_33 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  L0Memory_34 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  L0Memory_35 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  L0Memory_36 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  L0Memory_37 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  L0Memory_38 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  L0Memory_39 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  L0Memory_40 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  L0Memory_41 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  L0Memory_42 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  L0Memory_43 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  L0Memory_44 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  L0Memory_45 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  L0Memory_46 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  L0Memory_47 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  L0Memory_48 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  L0Memory_49 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  L0Memory_50 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  L0Memory_51 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  L0Memory_52 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  L0Memory_53 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  L0Memory_54 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  L0Memory_55 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  L0Memory_56 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  L0Memory_57 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  L0Memory_58 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  L0Memory_59 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  L0Memory_60 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  L0Memory_61 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  L0Memory_62 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  L0Memory_63 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  L0Memory_64 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  L0Memory_65 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  L0Memory_66 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  L0Memory_67 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  L0Memory_68 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  L0Memory_69 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  L0Memory_70 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  L0Memory_71 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  L0Memory_72 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  L0Memory_73 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  L0Memory_74 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  L0Memory_75 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  L0Memory_76 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  L0Memory_77 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  L0Memory_78 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  L0Memory_79 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  L0Memory_80 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  L0Memory_81 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  L0Memory_82 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  L0Memory_83 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  L0Memory_84 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  L0Memory_85 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  L0Memory_86 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  L0Memory_87 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  L0Memory_88 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  L0Memory_89 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  L0Memory_90 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  L0Memory_91 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  L0Memory_92 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  L0Memory_93 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  L0Memory_94 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  L0Memory_95 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  L0Memory_96 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  L0Memory_97 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  L0Memory_98 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  L0Memory_99 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  state = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  mux2out_reg = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  mux3out_reg = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  count = _RAND_104[9:0];
  _RAND_105 = {1{`RANDOM}};
  GRU_out_width = _RAND_105[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PE_2(
  input         clock,
  input         reset,
  input  [15:0] io_FromAbovePE,
  input  [15:0] io_FromL1,
  input  [2:0]  io_control_signal_control,
  input  [9:0]  io_control_signal_count,
  input  [5:0]  io_control_signal_L0index,
  input  [11:0] io_control_signal_mask,
  input  [7:0]  io_control_signal_gru_out_width,
  output [15:0] io_ToRightPE,
  output [15:0] io_ToBelowPE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] FP16MAC_io_a; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_b; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_c; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_out; // @[PEArray.scala 72:23]
  reg [5:0] L0Index; // @[PEArray.scala 39:24]
  reg [15:0] L0Memory_0; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_1; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_2; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_3; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_4; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_5; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_6; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_7; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_8; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_9; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_10; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_11; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_12; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_13; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_14; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_15; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_16; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_17; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_18; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_19; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_20; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_21; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_22; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_23; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_24; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_25; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_26; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_27; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_28; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_29; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_30; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_31; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_32; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_33; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_34; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_35; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_36; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_37; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_38; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_39; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_40; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_41; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_42; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_43; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_44; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_45; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_46; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_47; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_48; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_49; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_50; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_51; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_52; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_53; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_54; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_55; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_56; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_57; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_58; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_59; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_60; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_61; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_62; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_63; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_64; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_65; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_66; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_67; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_68; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_69; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_70; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_71; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_72; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_73; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_74; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_75; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_76; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_77; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_78; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_79; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_80; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_81; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_82; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_83; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_84; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_85; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_86; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_87; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_88; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_89; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_90; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_91; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_92; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_93; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_94; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_95; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_96; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_97; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_98; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_99; // @[PEArray.scala 40:21]
  reg [2:0] state; // @[PEArray.scala 100:22]
  wire  _T_3 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_12 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_16 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_22 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_31 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_41 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_342 = _T_41 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 231:12 PEArray.scala 32:8]
  wire  _GEN_349 = _T_31 ? 1'h0 : _GEN_342; // @[Conditional.scala 39:67 PEArray.scala 208:12]
  wire  _GEN_459 = _T_22 | _GEN_349; // @[Conditional.scala 39:67 PEArray.scala 32:8]
  wire  _GEN_572 = _T_12 | (_T_16 | _GEN_459); // @[Conditional.scala 39:67 PEArray.scala 149:12]
  wire  sel1 = _T_3 | _GEN_572; // @[Conditional.scala 40:58 PEArray.scala 108:12]
  wire [15:0] mux1out = sel1 ? io_FromL1 : 16'h0; // @[PEArray.scala 50:14 PEArray.scala 50:23 PEArray.scala 51:24]
  wire [15:0] MAC_out = FP16MAC_io_out; // @[PEArray.scala 47:21 PEArray.scala 85:11]
  wire  _GEN_465 = _T_16 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 177:12]
  wire  _GEN_580 = _T_12 | _GEN_465; // @[Conditional.scala 39:67 PEArray.scala 34:8]
  wire  sel3 = _T_3 | _GEN_580; // @[Conditional.scala 40:58 PEArray.scala 110:12]
  wire [1:0] _GEN_344 = _T_41 ? 2'h2 : 2'h0; // @[Conditional.scala 39:67 PEArray.scala 233:12 PEArray.scala 35:8]
  wire [1:0] _GEN_351 = _T_31 ? 2'h2 : _GEN_344; // @[Conditional.scala 39:67 PEArray.scala 210:12]
  wire [1:0] _GEN_461 = _T_22 ? 2'h0 : _GEN_351; // @[Conditional.scala 39:67 PEArray.scala 35:8]
  wire [1:0] _GEN_466 = _T_16 ? 2'h0 : _GEN_461; // @[Conditional.scala 39:67 PEArray.scala 178:12]
  wire [1:0] _GEN_574 = _T_12 ? 2'h1 : _GEN_466; // @[Conditional.scala 39:67]
  wire [1:0] sel4 = _T_3 ? 2'h0 : _GEN_574; // @[Conditional.scala 40:58 PEArray.scala 111:12]
  wire [15:0] _GEN_3 = sel4 == 2'h2 ? io_FromL1 : 16'h0; // @[PEArray.scala 65:28 PEArray.scala 66:15 PEArray.scala 69:15]
  wire [15:0] _GEN_4 = sel4 == 2'h1 ? io_FromAbovePE : _GEN_3; // @[PEArray.scala 62:28 PEArray.scala 63:15]
  wire [15:0] mux4out = sel4 == 2'h0 ? 16'h0 : _GEN_4; // @[PEArray.scala 59:22 PEArray.scala 60:13]
  wire [15:0] _GEN_7 = 6'h1 == L0Index ? L0Memory_1 : L0Memory_0; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_8 = 6'h2 == L0Index ? L0Memory_2 : _GEN_7; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_9 = 6'h3 == L0Index ? L0Memory_3 : _GEN_8; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_10 = 6'h4 == L0Index ? L0Memory_4 : _GEN_9; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_11 = 6'h5 == L0Index ? L0Memory_5 : _GEN_10; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_12 = 6'h6 == L0Index ? L0Memory_6 : _GEN_11; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_13 = 6'h7 == L0Index ? L0Memory_7 : _GEN_12; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_14 = 6'h8 == L0Index ? L0Memory_8 : _GEN_13; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_15 = 6'h9 == L0Index ? L0Memory_9 : _GEN_14; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_16 = 6'ha == L0Index ? L0Memory_10 : _GEN_15; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_17 = 6'hb == L0Index ? L0Memory_11 : _GEN_16; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_18 = 6'hc == L0Index ? L0Memory_12 : _GEN_17; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_19 = 6'hd == L0Index ? L0Memory_13 : _GEN_18; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_20 = 6'he == L0Index ? L0Memory_14 : _GEN_19; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_21 = 6'hf == L0Index ? L0Memory_15 : _GEN_20; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_22 = 6'h10 == L0Index ? L0Memory_16 : _GEN_21; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_23 = 6'h11 == L0Index ? L0Memory_17 : _GEN_22; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_24 = 6'h12 == L0Index ? L0Memory_18 : _GEN_23; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_25 = 6'h13 == L0Index ? L0Memory_19 : _GEN_24; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_26 = 6'h14 == L0Index ? L0Memory_20 : _GEN_25; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_27 = 6'h15 == L0Index ? L0Memory_21 : _GEN_26; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_28 = 6'h16 == L0Index ? L0Memory_22 : _GEN_27; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_29 = 6'h17 == L0Index ? L0Memory_23 : _GEN_28; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_30 = 6'h18 == L0Index ? L0Memory_24 : _GEN_29; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_31 = 6'h19 == L0Index ? L0Memory_25 : _GEN_30; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_32 = 6'h1a == L0Index ? L0Memory_26 : _GEN_31; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_33 = 6'h1b == L0Index ? L0Memory_27 : _GEN_32; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_34 = 6'h1c == L0Index ? L0Memory_28 : _GEN_33; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_35 = 6'h1d == L0Index ? L0Memory_29 : _GEN_34; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_36 = 6'h1e == L0Index ? L0Memory_30 : _GEN_35; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_37 = 6'h1f == L0Index ? L0Memory_31 : _GEN_36; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_38 = 6'h20 == L0Index ? L0Memory_32 : _GEN_37; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_39 = 6'h21 == L0Index ? L0Memory_33 : _GEN_38; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_40 = 6'h22 == L0Index ? L0Memory_34 : _GEN_39; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_41 = 6'h23 == L0Index ? L0Memory_35 : _GEN_40; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_42 = 6'h24 == L0Index ? L0Memory_36 : _GEN_41; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_43 = 6'h25 == L0Index ? L0Memory_37 : _GEN_42; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_44 = 6'h26 == L0Index ? L0Memory_38 : _GEN_43; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_45 = 6'h27 == L0Index ? L0Memory_39 : _GEN_44; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_46 = 6'h28 == L0Index ? L0Memory_40 : _GEN_45; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_47 = 6'h29 == L0Index ? L0Memory_41 : _GEN_46; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_48 = 6'h2a == L0Index ? L0Memory_42 : _GEN_47; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_49 = 6'h2b == L0Index ? L0Memory_43 : _GEN_48; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_50 = 6'h2c == L0Index ? L0Memory_44 : _GEN_49; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_51 = 6'h2d == L0Index ? L0Memory_45 : _GEN_50; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_52 = 6'h2e == L0Index ? L0Memory_46 : _GEN_51; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_53 = 6'h2f == L0Index ? L0Memory_47 : _GEN_52; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_54 = 6'h30 == L0Index ? L0Memory_48 : _GEN_53; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_55 = 6'h31 == L0Index ? L0Memory_49 : _GEN_54; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_56 = 6'h32 == L0Index ? L0Memory_50 : _GEN_55; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_57 = 6'h33 == L0Index ? L0Memory_51 : _GEN_56; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_58 = 6'h34 == L0Index ? L0Memory_52 : _GEN_57; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_59 = 6'h35 == L0Index ? L0Memory_53 : _GEN_58; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_60 = 6'h36 == L0Index ? L0Memory_54 : _GEN_59; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_61 = 6'h37 == L0Index ? L0Memory_55 : _GEN_60; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_62 = 6'h38 == L0Index ? L0Memory_56 : _GEN_61; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_63 = 6'h39 == L0Index ? L0Memory_57 : _GEN_62; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_64 = 6'h3a == L0Index ? L0Memory_58 : _GEN_63; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_65 = 6'h3b == L0Index ? L0Memory_59 : _GEN_64; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_66 = 6'h3c == L0Index ? L0Memory_60 : _GEN_65; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_67 = 6'h3d == L0Index ? L0Memory_61 : _GEN_66; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_68 = 6'h3e == L0Index ? L0Memory_62 : _GEN_67; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_69 = 6'h3f == L0Index ? L0Memory_63 : _GEN_68; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [6:0] _GEN_793 = {{1'd0}, L0Index}; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_70 = 7'h40 == _GEN_793 ? L0Memory_64 : _GEN_69; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_71 = 7'h41 == _GEN_793 ? L0Memory_65 : _GEN_70; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_72 = 7'h42 == _GEN_793 ? L0Memory_66 : _GEN_71; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_73 = 7'h43 == _GEN_793 ? L0Memory_67 : _GEN_72; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_74 = 7'h44 == _GEN_793 ? L0Memory_68 : _GEN_73; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_75 = 7'h45 == _GEN_793 ? L0Memory_69 : _GEN_74; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_76 = 7'h46 == _GEN_793 ? L0Memory_70 : _GEN_75; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_77 = 7'h47 == _GEN_793 ? L0Memory_71 : _GEN_76; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_78 = 7'h48 == _GEN_793 ? L0Memory_72 : _GEN_77; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_79 = 7'h49 == _GEN_793 ? L0Memory_73 : _GEN_78; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_80 = 7'h4a == _GEN_793 ? L0Memory_74 : _GEN_79; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_81 = 7'h4b == _GEN_793 ? L0Memory_75 : _GEN_80; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_82 = 7'h4c == _GEN_793 ? L0Memory_76 : _GEN_81; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_83 = 7'h4d == _GEN_793 ? L0Memory_77 : _GEN_82; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_84 = 7'h4e == _GEN_793 ? L0Memory_78 : _GEN_83; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_85 = 7'h4f == _GEN_793 ? L0Memory_79 : _GEN_84; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_86 = 7'h50 == _GEN_793 ? L0Memory_80 : _GEN_85; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_87 = 7'h51 == _GEN_793 ? L0Memory_81 : _GEN_86; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_88 = 7'h52 == _GEN_793 ? L0Memory_82 : _GEN_87; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_89 = 7'h53 == _GEN_793 ? L0Memory_83 : _GEN_88; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_90 = 7'h54 == _GEN_793 ? L0Memory_84 : _GEN_89; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_91 = 7'h55 == _GEN_793 ? L0Memory_85 : _GEN_90; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_92 = 7'h56 == _GEN_793 ? L0Memory_86 : _GEN_91; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_93 = 7'h57 == _GEN_793 ? L0Memory_87 : _GEN_92; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_94 = 7'h58 == _GEN_793 ? L0Memory_88 : _GEN_93; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_95 = 7'h59 == _GEN_793 ? L0Memory_89 : _GEN_94; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_96 = 7'h5a == _GEN_793 ? L0Memory_90 : _GEN_95; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_97 = 7'h5b == _GEN_793 ? L0Memory_91 : _GEN_96; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_98 = 7'h5c == _GEN_793 ? L0Memory_92 : _GEN_97; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_99 = 7'h5d == _GEN_793 ? L0Memory_93 : _GEN_98; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_100 = 7'h5e == _GEN_793 ? L0Memory_94 : _GEN_99; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_101 = 7'h5f == _GEN_793 ? L0Memory_95 : _GEN_100; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_102 = 7'h60 == _GEN_793 ? L0Memory_96 : _GEN_101; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_103 = 7'h61 == _GEN_793 ? L0Memory_97 : _GEN_102; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_104 = 7'h62 == _GEN_793 ? L0Memory_98 : _GEN_103; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_105 = 7'h63 == _GEN_793 ? L0Memory_99 : _GEN_104; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire  _GEN_467 = _T_16 ? 1'h0 : _GEN_459; // @[Conditional.scala 39:67 PEArray.scala 179:12]
  wire  _GEN_575 = _T_12 ? 1'h0 : _GEN_467; // @[Conditional.scala 39:67 PEArray.scala 157:12]
  wire  sel5 = _T_3 ? 1'h0 : _GEN_575; // @[Conditional.scala 40:58 PEArray.scala 112:12]
  reg [15:0] mux2out_reg; // @[PEArray.scala 90:28]
  reg [15:0] mux3out_reg; // @[PEArray.scala 91:28]
  reg [9:0] count; // @[PEArray.scala 101:22]
  reg [9:0] count_max; // @[PEArray.scala 102:22]
  reg [5:0] L0index_begin; // @[PEArray.scala 103:26]
  reg [5:0] GRU_out_width; // @[PEArray.scala 104:26]
  wire  _T_6 = 3'h0 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_7 = 3'h1 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_8 = 3'h2 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_9 = 3'h3 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_10 = 3'h4 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_11 = 3'h5 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_109 = _T_11 ? 3'h5 : state; // @[Conditional.scala 39:67 PEArray.scala 140:19 PEArray.scala 100:22]
  wire [2:0] _GEN_110 = _T_10 ? 3'h4 : _GEN_109; // @[Conditional.scala 39:67 PEArray.scala 136:19]
  wire [2:0] _GEN_111 = _T_9 ? 3'h3 : _GEN_110; // @[Conditional.scala 39:67 PEArray.scala 132:19]
  wire [2:0] _GEN_112 = _T_8 ? 3'h2 : _GEN_111; // @[Conditional.scala 39:67 PEArray.scala 128:19]
  wire [2:0] _GEN_113 = _T_7 ? 3'h1 : _GEN_112; // @[Conditional.scala 39:67 PEArray.scala 124:19]
  wire [7:0] _GEN_118 = io_control_signal_mask[11] ? io_control_signal_gru_out_width : {{2'd0}, GRU_out_width}; // @[PEArray.scala 116:57 PEArray.scala 145:23 PEArray.scala 104:26]
  wire [9:0] _count_T_1 = count + 10'h1; // @[PEArray.scala 162:24]
  wire [9:0] _GEN_120 = count != 10'h33 ? _count_T_1 : count; // @[PEArray.scala 161:27 PEArray.scala 162:15 PEArray.scala 101:22]
  wire [9:0] _GEN_124 = count != 10'h188 ? _count_T_1 : count; // @[PEArray.scala 183:28 PEArray.scala 184:15 PEArray.scala 101:22]
  wire [9:0] _GEN_125 = count == 10'h188 ? 10'h0 : _GEN_124; // @[PEArray.scala 186:28 PEArray.scala 187:15]
  wire [2:0] _GEN_126 = count == 10'h188 ? 3'h0 : state; // @[PEArray.scala 186:28 PEArray.scala 188:15 PEArray.scala 100:22]
  wire [9:0] _GEN_127 = count != count_max ? _count_T_1 : count; // @[PEArray.scala 192:32 PEArray.scala 193:15 PEArray.scala 101:22]
  wire [5:0] _GEN_128 = count == 10'h0 ? L0index_begin : L0Index; // @[PEArray.scala 195:26 PEArray.scala 196:17 PEArray.scala 39:24]
  wire [9:0] _T_27 = count_max - 10'h1; // @[PEArray.scala 198:51]
  wire [15:0] _GEN_129 = 6'h0 == L0Index ? io_FromL1 : L0Memory_0; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_130 = 6'h1 == L0Index ? io_FromL1 : L0Memory_1; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_131 = 6'h2 == L0Index ? io_FromL1 : L0Memory_2; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_132 = 6'h3 == L0Index ? io_FromL1 : L0Memory_3; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_133 = 6'h4 == L0Index ? io_FromL1 : L0Memory_4; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_134 = 6'h5 == L0Index ? io_FromL1 : L0Memory_5; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_135 = 6'h6 == L0Index ? io_FromL1 : L0Memory_6; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_136 = 6'h7 == L0Index ? io_FromL1 : L0Memory_7; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_137 = 6'h8 == L0Index ? io_FromL1 : L0Memory_8; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_138 = 6'h9 == L0Index ? io_FromL1 : L0Memory_9; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_139 = 6'ha == L0Index ? io_FromL1 : L0Memory_10; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_140 = 6'hb == L0Index ? io_FromL1 : L0Memory_11; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_141 = 6'hc == L0Index ? io_FromL1 : L0Memory_12; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_142 = 6'hd == L0Index ? io_FromL1 : L0Memory_13; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_143 = 6'he == L0Index ? io_FromL1 : L0Memory_14; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_144 = 6'hf == L0Index ? io_FromL1 : L0Memory_15; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_145 = 6'h10 == L0Index ? io_FromL1 : L0Memory_16; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_146 = 6'h11 == L0Index ? io_FromL1 : L0Memory_17; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_147 = 6'h12 == L0Index ? io_FromL1 : L0Memory_18; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_148 = 6'h13 == L0Index ? io_FromL1 : L0Memory_19; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_149 = 6'h14 == L0Index ? io_FromL1 : L0Memory_20; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_150 = 6'h15 == L0Index ? io_FromL1 : L0Memory_21; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_151 = 6'h16 == L0Index ? io_FromL1 : L0Memory_22; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_152 = 6'h17 == L0Index ? io_FromL1 : L0Memory_23; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_153 = 6'h18 == L0Index ? io_FromL1 : L0Memory_24; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_154 = 6'h19 == L0Index ? io_FromL1 : L0Memory_25; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_155 = 6'h1a == L0Index ? io_FromL1 : L0Memory_26; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_156 = 6'h1b == L0Index ? io_FromL1 : L0Memory_27; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_157 = 6'h1c == L0Index ? io_FromL1 : L0Memory_28; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_158 = 6'h1d == L0Index ? io_FromL1 : L0Memory_29; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_159 = 6'h1e == L0Index ? io_FromL1 : L0Memory_30; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_160 = 6'h1f == L0Index ? io_FromL1 : L0Memory_31; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_161 = 6'h20 == L0Index ? io_FromL1 : L0Memory_32; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_162 = 6'h21 == L0Index ? io_FromL1 : L0Memory_33; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_163 = 6'h22 == L0Index ? io_FromL1 : L0Memory_34; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_164 = 6'h23 == L0Index ? io_FromL1 : L0Memory_35; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_165 = 6'h24 == L0Index ? io_FromL1 : L0Memory_36; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_166 = 6'h25 == L0Index ? io_FromL1 : L0Memory_37; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_167 = 6'h26 == L0Index ? io_FromL1 : L0Memory_38; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_168 = 6'h27 == L0Index ? io_FromL1 : L0Memory_39; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_169 = 6'h28 == L0Index ? io_FromL1 : L0Memory_40; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_170 = 6'h29 == L0Index ? io_FromL1 : L0Memory_41; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_171 = 6'h2a == L0Index ? io_FromL1 : L0Memory_42; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_172 = 6'h2b == L0Index ? io_FromL1 : L0Memory_43; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_173 = 6'h2c == L0Index ? io_FromL1 : L0Memory_44; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_174 = 6'h2d == L0Index ? io_FromL1 : L0Memory_45; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_175 = 6'h2e == L0Index ? io_FromL1 : L0Memory_46; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_176 = 6'h2f == L0Index ? io_FromL1 : L0Memory_47; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_177 = 6'h30 == L0Index ? io_FromL1 : L0Memory_48; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_178 = 6'h31 == L0Index ? io_FromL1 : L0Memory_49; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_179 = 6'h32 == L0Index ? io_FromL1 : L0Memory_50; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_180 = 6'h33 == L0Index ? io_FromL1 : L0Memory_51; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_181 = 6'h34 == L0Index ? io_FromL1 : L0Memory_52; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_182 = 6'h35 == L0Index ? io_FromL1 : L0Memory_53; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_183 = 6'h36 == L0Index ? io_FromL1 : L0Memory_54; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_184 = 6'h37 == L0Index ? io_FromL1 : L0Memory_55; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_185 = 6'h38 == L0Index ? io_FromL1 : L0Memory_56; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_186 = 6'h39 == L0Index ? io_FromL1 : L0Memory_57; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_187 = 6'h3a == L0Index ? io_FromL1 : L0Memory_58; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_188 = 6'h3b == L0Index ? io_FromL1 : L0Memory_59; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_189 = 6'h3c == L0Index ? io_FromL1 : L0Memory_60; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_190 = 6'h3d == L0Index ? io_FromL1 : L0Memory_61; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_191 = 6'h3e == L0Index ? io_FromL1 : L0Memory_62; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_192 = 6'h3f == L0Index ? io_FromL1 : L0Memory_63; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_193 = 7'h40 == _GEN_793 ? io_FromL1 : L0Memory_64; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_194 = 7'h41 == _GEN_793 ? io_FromL1 : L0Memory_65; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_195 = 7'h42 == _GEN_793 ? io_FromL1 : L0Memory_66; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_196 = 7'h43 == _GEN_793 ? io_FromL1 : L0Memory_67; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_197 = 7'h44 == _GEN_793 ? io_FromL1 : L0Memory_68; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_198 = 7'h45 == _GEN_793 ? io_FromL1 : L0Memory_69; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_199 = 7'h46 == _GEN_793 ? io_FromL1 : L0Memory_70; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_200 = 7'h47 == _GEN_793 ? io_FromL1 : L0Memory_71; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_201 = 7'h48 == _GEN_793 ? io_FromL1 : L0Memory_72; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_202 = 7'h49 == _GEN_793 ? io_FromL1 : L0Memory_73; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_203 = 7'h4a == _GEN_793 ? io_FromL1 : L0Memory_74; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_204 = 7'h4b == _GEN_793 ? io_FromL1 : L0Memory_75; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_205 = 7'h4c == _GEN_793 ? io_FromL1 : L0Memory_76; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_206 = 7'h4d == _GEN_793 ? io_FromL1 : L0Memory_77; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_207 = 7'h4e == _GEN_793 ? io_FromL1 : L0Memory_78; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_208 = 7'h4f == _GEN_793 ? io_FromL1 : L0Memory_79; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_209 = 7'h50 == _GEN_793 ? io_FromL1 : L0Memory_80; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_210 = 7'h51 == _GEN_793 ? io_FromL1 : L0Memory_81; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_211 = 7'h52 == _GEN_793 ? io_FromL1 : L0Memory_82; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_212 = 7'h53 == _GEN_793 ? io_FromL1 : L0Memory_83; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_213 = 7'h54 == _GEN_793 ? io_FromL1 : L0Memory_84; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_214 = 7'h55 == _GEN_793 ? io_FromL1 : L0Memory_85; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_215 = 7'h56 == _GEN_793 ? io_FromL1 : L0Memory_86; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_216 = 7'h57 == _GEN_793 ? io_FromL1 : L0Memory_87; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_217 = 7'h58 == _GEN_793 ? io_FromL1 : L0Memory_88; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_218 = 7'h59 == _GEN_793 ? io_FromL1 : L0Memory_89; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_219 = 7'h5a == _GEN_793 ? io_FromL1 : L0Memory_90; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_220 = 7'h5b == _GEN_793 ? io_FromL1 : L0Memory_91; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_221 = 7'h5c == _GEN_793 ? io_FromL1 : L0Memory_92; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_222 = 7'h5d == _GEN_793 ? io_FromL1 : L0Memory_93; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_223 = 7'h5e == _GEN_793 ? io_FromL1 : L0Memory_94; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_224 = 7'h5f == _GEN_793 ? io_FromL1 : L0Memory_95; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_225 = 7'h60 == _GEN_793 ? io_FromL1 : L0Memory_96; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_226 = 7'h61 == _GEN_793 ? io_FromL1 : L0Memory_97; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_227 = 7'h62 == _GEN_793 ? io_FromL1 : L0Memory_98; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_228 = 7'h63 == _GEN_793 ? io_FromL1 : L0Memory_99; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [5:0] _L0Index_T_2 = L0Index + 6'h1; // @[PEArray.scala 200:28]
  wire [15:0] _GEN_229 = count >= 10'h1 & count <= _T_27 ? _GEN_129 : L0Memory_0; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_230 = count >= 10'h1 & count <= _T_27 ? _GEN_130 : L0Memory_1; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_231 = count >= 10'h1 & count <= _T_27 ? _GEN_131 : L0Memory_2; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_232 = count >= 10'h1 & count <= _T_27 ? _GEN_132 : L0Memory_3; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_233 = count >= 10'h1 & count <= _T_27 ? _GEN_133 : L0Memory_4; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_234 = count >= 10'h1 & count <= _T_27 ? _GEN_134 : L0Memory_5; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_235 = count >= 10'h1 & count <= _T_27 ? _GEN_135 : L0Memory_6; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_236 = count >= 10'h1 & count <= _T_27 ? _GEN_136 : L0Memory_7; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_237 = count >= 10'h1 & count <= _T_27 ? _GEN_137 : L0Memory_8; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_238 = count >= 10'h1 & count <= _T_27 ? _GEN_138 : L0Memory_9; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_239 = count >= 10'h1 & count <= _T_27 ? _GEN_139 : L0Memory_10; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_240 = count >= 10'h1 & count <= _T_27 ? _GEN_140 : L0Memory_11; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_241 = count >= 10'h1 & count <= _T_27 ? _GEN_141 : L0Memory_12; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_242 = count >= 10'h1 & count <= _T_27 ? _GEN_142 : L0Memory_13; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_243 = count >= 10'h1 & count <= _T_27 ? _GEN_143 : L0Memory_14; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_244 = count >= 10'h1 & count <= _T_27 ? _GEN_144 : L0Memory_15; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_245 = count >= 10'h1 & count <= _T_27 ? _GEN_145 : L0Memory_16; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_246 = count >= 10'h1 & count <= _T_27 ? _GEN_146 : L0Memory_17; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_247 = count >= 10'h1 & count <= _T_27 ? _GEN_147 : L0Memory_18; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_248 = count >= 10'h1 & count <= _T_27 ? _GEN_148 : L0Memory_19; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_249 = count >= 10'h1 & count <= _T_27 ? _GEN_149 : L0Memory_20; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_250 = count >= 10'h1 & count <= _T_27 ? _GEN_150 : L0Memory_21; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_251 = count >= 10'h1 & count <= _T_27 ? _GEN_151 : L0Memory_22; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_252 = count >= 10'h1 & count <= _T_27 ? _GEN_152 : L0Memory_23; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_253 = count >= 10'h1 & count <= _T_27 ? _GEN_153 : L0Memory_24; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_254 = count >= 10'h1 & count <= _T_27 ? _GEN_154 : L0Memory_25; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_255 = count >= 10'h1 & count <= _T_27 ? _GEN_155 : L0Memory_26; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_256 = count >= 10'h1 & count <= _T_27 ? _GEN_156 : L0Memory_27; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_257 = count >= 10'h1 & count <= _T_27 ? _GEN_157 : L0Memory_28; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_258 = count >= 10'h1 & count <= _T_27 ? _GEN_158 : L0Memory_29; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_259 = count >= 10'h1 & count <= _T_27 ? _GEN_159 : L0Memory_30; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_260 = count >= 10'h1 & count <= _T_27 ? _GEN_160 : L0Memory_31; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_261 = count >= 10'h1 & count <= _T_27 ? _GEN_161 : L0Memory_32; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_262 = count >= 10'h1 & count <= _T_27 ? _GEN_162 : L0Memory_33; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_263 = count >= 10'h1 & count <= _T_27 ? _GEN_163 : L0Memory_34; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_264 = count >= 10'h1 & count <= _T_27 ? _GEN_164 : L0Memory_35; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_265 = count >= 10'h1 & count <= _T_27 ? _GEN_165 : L0Memory_36; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_266 = count >= 10'h1 & count <= _T_27 ? _GEN_166 : L0Memory_37; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_267 = count >= 10'h1 & count <= _T_27 ? _GEN_167 : L0Memory_38; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_268 = count >= 10'h1 & count <= _T_27 ? _GEN_168 : L0Memory_39; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_269 = count >= 10'h1 & count <= _T_27 ? _GEN_169 : L0Memory_40; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_270 = count >= 10'h1 & count <= _T_27 ? _GEN_170 : L0Memory_41; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_271 = count >= 10'h1 & count <= _T_27 ? _GEN_171 : L0Memory_42; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_272 = count >= 10'h1 & count <= _T_27 ? _GEN_172 : L0Memory_43; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_273 = count >= 10'h1 & count <= _T_27 ? _GEN_173 : L0Memory_44; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_274 = count >= 10'h1 & count <= _T_27 ? _GEN_174 : L0Memory_45; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_275 = count >= 10'h1 & count <= _T_27 ? _GEN_175 : L0Memory_46; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_276 = count >= 10'h1 & count <= _T_27 ? _GEN_176 : L0Memory_47; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_277 = count >= 10'h1 & count <= _T_27 ? _GEN_177 : L0Memory_48; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_278 = count >= 10'h1 & count <= _T_27 ? _GEN_178 : L0Memory_49; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_279 = count >= 10'h1 & count <= _T_27 ? _GEN_179 : L0Memory_50; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_280 = count >= 10'h1 & count <= _T_27 ? _GEN_180 : L0Memory_51; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_281 = count >= 10'h1 & count <= _T_27 ? _GEN_181 : L0Memory_52; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_282 = count >= 10'h1 & count <= _T_27 ? _GEN_182 : L0Memory_53; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_283 = count >= 10'h1 & count <= _T_27 ? _GEN_183 : L0Memory_54; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_284 = count >= 10'h1 & count <= _T_27 ? _GEN_184 : L0Memory_55; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_285 = count >= 10'h1 & count <= _T_27 ? _GEN_185 : L0Memory_56; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_286 = count >= 10'h1 & count <= _T_27 ? _GEN_186 : L0Memory_57; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_287 = count >= 10'h1 & count <= _T_27 ? _GEN_187 : L0Memory_58; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_288 = count >= 10'h1 & count <= _T_27 ? _GEN_188 : L0Memory_59; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_289 = count >= 10'h1 & count <= _T_27 ? _GEN_189 : L0Memory_60; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_290 = count >= 10'h1 & count <= _T_27 ? _GEN_190 : L0Memory_61; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_291 = count >= 10'h1 & count <= _T_27 ? _GEN_191 : L0Memory_62; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_292 = count >= 10'h1 & count <= _T_27 ? _GEN_192 : L0Memory_63; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_293 = count >= 10'h1 & count <= _T_27 ? _GEN_193 : L0Memory_64; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_294 = count >= 10'h1 & count <= _T_27 ? _GEN_194 : L0Memory_65; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_295 = count >= 10'h1 & count <= _T_27 ? _GEN_195 : L0Memory_66; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_296 = count >= 10'h1 & count <= _T_27 ? _GEN_196 : L0Memory_67; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_297 = count >= 10'h1 & count <= _T_27 ? _GEN_197 : L0Memory_68; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_298 = count >= 10'h1 & count <= _T_27 ? _GEN_198 : L0Memory_69; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_299 = count >= 10'h1 & count <= _T_27 ? _GEN_199 : L0Memory_70; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_300 = count >= 10'h1 & count <= _T_27 ? _GEN_200 : L0Memory_71; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_301 = count >= 10'h1 & count <= _T_27 ? _GEN_201 : L0Memory_72; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_302 = count >= 10'h1 & count <= _T_27 ? _GEN_202 : L0Memory_73; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_303 = count >= 10'h1 & count <= _T_27 ? _GEN_203 : L0Memory_74; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_304 = count >= 10'h1 & count <= _T_27 ? _GEN_204 : L0Memory_75; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_305 = count >= 10'h1 & count <= _T_27 ? _GEN_205 : L0Memory_76; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_306 = count >= 10'h1 & count <= _T_27 ? _GEN_206 : L0Memory_77; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_307 = count >= 10'h1 & count <= _T_27 ? _GEN_207 : L0Memory_78; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_308 = count >= 10'h1 & count <= _T_27 ? _GEN_208 : L0Memory_79; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_309 = count >= 10'h1 & count <= _T_27 ? _GEN_209 : L0Memory_80; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_310 = count >= 10'h1 & count <= _T_27 ? _GEN_210 : L0Memory_81; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_311 = count >= 10'h1 & count <= _T_27 ? _GEN_211 : L0Memory_82; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_312 = count >= 10'h1 & count <= _T_27 ? _GEN_212 : L0Memory_83; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_313 = count >= 10'h1 & count <= _T_27 ? _GEN_213 : L0Memory_84; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_314 = count >= 10'h1 & count <= _T_27 ? _GEN_214 : L0Memory_85; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_315 = count >= 10'h1 & count <= _T_27 ? _GEN_215 : L0Memory_86; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_316 = count >= 10'h1 & count <= _T_27 ? _GEN_216 : L0Memory_87; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_317 = count >= 10'h1 & count <= _T_27 ? _GEN_217 : L0Memory_88; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_318 = count >= 10'h1 & count <= _T_27 ? _GEN_218 : L0Memory_89; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_319 = count >= 10'h1 & count <= _T_27 ? _GEN_219 : L0Memory_90; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_320 = count >= 10'h1 & count <= _T_27 ? _GEN_220 : L0Memory_91; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_321 = count >= 10'h1 & count <= _T_27 ? _GEN_221 : L0Memory_92; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_322 = count >= 10'h1 & count <= _T_27 ? _GEN_222 : L0Memory_93; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_323 = count >= 10'h1 & count <= _T_27 ? _GEN_223 : L0Memory_94; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_324 = count >= 10'h1 & count <= _T_27 ? _GEN_224 : L0Memory_95; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_325 = count >= 10'h1 & count <= _T_27 ? _GEN_225 : L0Memory_96; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_326 = count >= 10'h1 & count <= _T_27 ? _GEN_226 : L0Memory_97; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_327 = count >= 10'h1 & count <= _T_27 ? _GEN_227 : L0Memory_98; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_328 = count >= 10'h1 & count <= _T_27 ? _GEN_228 : L0Memory_99; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [5:0] _GEN_329 = count >= 10'h1 & count <= _T_27 ? _L0Index_T_2 : _GEN_128; // @[PEArray.scala 198:59 PEArray.scala 200:17]
  wire [9:0] _GEN_330 = count == count_max ? 10'h0 : _GEN_127; // @[PEArray.scala 202:32 PEArray.scala 203:15]
  wire [2:0] _GEN_331 = count == count_max ? 3'h0 : state; // @[PEArray.scala 202:32 PEArray.scala 204:15 PEArray.scala 100:22]
  wire [9:0] _GEN_865 = {{4'd0}, GRU_out_width}; // @[PEArray.scala 220:19]
  wire [9:0] _GEN_0 = count % _GEN_865; // @[PEArray.scala 220:19]
  wire [5:0] _T_36 = _GEN_0[5:0]; // @[PEArray.scala 220:19]
  wire [5:0] _T_38 = GRU_out_width - 6'h1; // @[PEArray.scala 220:55]
  wire [5:0] _GEN_334 = _T_36 == _T_38 ? _L0Index_T_2 : L0index_begin; // @[PEArray.scala 220:62 PEArray.scala 221:17 PEArray.scala 214:15]
  wire [5:0] _GEN_346 = _T_41 ? _GEN_334 : L0Index; // @[Conditional.scala 39:67 PEArray.scala 39:24]
  wire [9:0] _GEN_347 = _T_41 ? _GEN_330 : count; // @[Conditional.scala 39:67 PEArray.scala 101:22]
  wire [2:0] _GEN_348 = _T_41 ? _GEN_331 : state; // @[Conditional.scala 39:67 PEArray.scala 100:22]
  wire [5:0] _GEN_353 = _T_31 ? _GEN_334 : _GEN_346; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_354 = _T_31 ? _GEN_330 : _GEN_347; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_355 = _T_31 ? _GEN_331 : _GEN_348; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_356 = _T_22 ? _GEN_330 : _GEN_354; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_357 = _T_22 ? _GEN_329 : _GEN_353; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_458 = _T_22 ? _GEN_331 : _GEN_355; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_690 = _T_3 ? _GEN_118 : {{2'd0}, GRU_out_width}; // @[Conditional.scala 40:58 PEArray.scala 104:26]
  FP16MulAdder FP16MAC ( // @[PEArray.scala 72:23]
    .io_a(FP16MAC_io_a),
    .io_b(FP16MAC_io_b),
    .io_c(FP16MAC_io_c),
    .io_out(FP16MAC_io_out)
  );
  assign io_ToRightPE = mux3out_reg; // @[PEArray.scala 95:16]
  assign io_ToBelowPE = mux2out_reg; // @[PEArray.scala 94:16]
  assign FP16MAC_io_a = sel1 ? mux1out : 16'h0; // @[PEArray.scala 87:14 PEArray.scala 87:23 PEArray.scala 88:24]
  assign FP16MAC_io_b = sel5 ? mux4out : _GEN_105; // @[PEArray.scala 77:13 PEArray.scala 78:18 PEArray.scala 81:18]
  assign FP16MAC_io_c = sel5 ? _GEN_105 : mux4out; // @[PEArray.scala 77:13 PEArray.scala 79:18 PEArray.scala 82:18]
  always @(posedge clock) begin
    if (reset) begin // @[PEArray.scala 39:24]
      L0Index <= 6'h0; // @[PEArray.scala 39:24]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h2; // @[PEArray.scala 159:15]
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h3; // @[PEArray.scala 181:15]
      end else begin
        L0Index <= _GEN_357;
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_0 <= _GEN_229;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_1 <= _GEN_230;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_2 <= _GEN_231;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_3 <= _GEN_232;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_4 <= _GEN_233;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_5 <= _GEN_234;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_6 <= _GEN_235;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_7 <= _GEN_236;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_8 <= _GEN_237;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_9 <= _GEN_238;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_10 <= _GEN_239;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_11 <= _GEN_240;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_12 <= _GEN_241;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_13 <= _GEN_242;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_14 <= _GEN_243;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_15 <= _GEN_244;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_16 <= _GEN_245;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_17 <= _GEN_246;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_18 <= _GEN_247;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_19 <= _GEN_248;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_20 <= _GEN_249;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_21 <= _GEN_250;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_22 <= _GEN_251;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_23 <= _GEN_252;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_24 <= _GEN_253;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_25 <= _GEN_254;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_26 <= _GEN_255;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_27 <= _GEN_256;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_28 <= _GEN_257;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_29 <= _GEN_258;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_30 <= _GEN_259;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_31 <= _GEN_260;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_32 <= _GEN_261;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_33 <= _GEN_262;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_34 <= _GEN_263;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_35 <= _GEN_264;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_36 <= _GEN_265;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_37 <= _GEN_266;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_38 <= _GEN_267;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_39 <= _GEN_268;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_40 <= _GEN_269;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_41 <= _GEN_270;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_42 <= _GEN_271;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_43 <= _GEN_272;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_44 <= _GEN_273;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_45 <= _GEN_274;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_46 <= _GEN_275;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_47 <= _GEN_276;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_48 <= _GEN_277;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_49 <= _GEN_278;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_50 <= _GEN_279;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_51 <= _GEN_280;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_52 <= _GEN_281;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_53 <= _GEN_282;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_54 <= _GEN_283;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_55 <= _GEN_284;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_56 <= _GEN_285;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_57 <= _GEN_286;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_58 <= _GEN_287;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_59 <= _GEN_288;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_60 <= _GEN_289;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_61 <= _GEN_290;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_62 <= _GEN_291;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_63 <= _GEN_292;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_64 <= _GEN_293;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_65 <= _GEN_294;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_66 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_67 <= _GEN_296;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_68 <= _GEN_297;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_69 <= _GEN_298;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_70 <= _GEN_299;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_71 <= _GEN_300;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_72 <= _GEN_301;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_73 <= _GEN_302;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_74 <= _GEN_303;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_75 <= _GEN_304;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_76 <= _GEN_305;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_77 <= _GEN_306;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_78 <= _GEN_307;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_79 <= _GEN_308;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_80 <= _GEN_309;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_81 <= _GEN_310;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_82 <= _GEN_311;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_83 <= _GEN_312;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_84 <= _GEN_313;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_85 <= _GEN_314;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_86 <= _GEN_315;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_87 <= _GEN_316;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_88 <= _GEN_317;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_89 <= _GEN_318;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_90 <= _GEN_319;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_91 <= _GEN_320;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_92 <= _GEN_321;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_93 <= _GEN_322;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_94 <= _GEN_323;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_95 <= _GEN_324;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_96 <= _GEN_325;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_97 <= _GEN_326;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_98 <= _GEN_327;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_99 <= _GEN_328;
          end
        end
      end
    end
    if (reset) begin // @[PEArray.scala 100:22]
      state <= 3'h0; // @[PEArray.scala 100:22]
    end else if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[11]) begin // @[PEArray.scala 116:57]
        if (_T_6) begin // @[Conditional.scala 40:58]
          state <= 3'h0; // @[PEArray.scala 120:19]
        end else begin
          state <= _GEN_113;
        end
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      if (count == 10'h33) begin // @[PEArray.scala 164:27]
        state <= 3'h0; // @[PEArray.scala 166:15]
      end
    end else if (_T_16) begin // @[Conditional.scala 39:67]
      state <= _GEN_126;
    end else begin
      state <= _GEN_458;
    end
    if (reset) begin // @[PEArray.scala 90:28]
      mux2out_reg <= 16'h0; // @[PEArray.scala 90:28]
    end else begin
      mux2out_reg <= MAC_out; // @[PEArray.scala 90:28]
    end
    if (reset) begin // @[PEArray.scala 91:28]
      mux3out_reg <= 16'h0; // @[PEArray.scala 91:28]
    end else if (sel3) begin // @[PEArray.scala 56:14]
      mux3out_reg <= MAC_out; // @[PEArray.scala 56:23]
    end else if (sel1) begin // @[PEArray.scala 50:14]
      mux3out_reg <= io_FromL1; // @[PEArray.scala 50:23]
    end else begin
      mux3out_reg <= 16'h0; // @[PEArray.scala 51:24]
    end
    if (reset) begin // @[PEArray.scala 101:22]
      count <= 10'h0; // @[PEArray.scala 101:22]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        if (count == 10'h33) begin // @[PEArray.scala 164:27]
          count <= 10'h0; // @[PEArray.scala 165:15]
        end else begin
          count <= _GEN_120;
        end
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        count <= _GEN_125;
      end else begin
        count <= _GEN_356;
      end
    end
    if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[11]) begin // @[PEArray.scala 116:57]
        count_max <= io_control_signal_count; // @[PEArray.scala 143:19]
      end
    end
    if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[11]) begin // @[PEArray.scala 116:57]
        L0index_begin <= io_control_signal_L0index; // @[PEArray.scala 144:23]
      end
    end
    GRU_out_width <= _GEN_690[5:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  L0Index = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  L0Memory_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  L0Memory_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  L0Memory_2 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  L0Memory_3 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  L0Memory_4 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  L0Memory_5 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  L0Memory_6 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  L0Memory_7 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  L0Memory_8 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  L0Memory_9 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  L0Memory_10 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  L0Memory_11 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  L0Memory_12 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  L0Memory_13 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  L0Memory_14 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  L0Memory_15 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  L0Memory_16 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  L0Memory_17 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  L0Memory_18 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  L0Memory_19 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  L0Memory_20 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  L0Memory_21 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  L0Memory_22 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  L0Memory_23 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  L0Memory_24 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  L0Memory_25 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  L0Memory_26 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  L0Memory_27 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  L0Memory_28 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  L0Memory_29 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  L0Memory_30 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  L0Memory_31 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  L0Memory_32 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  L0Memory_33 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  L0Memory_34 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  L0Memory_35 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  L0Memory_36 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  L0Memory_37 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  L0Memory_38 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  L0Memory_39 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  L0Memory_40 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  L0Memory_41 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  L0Memory_42 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  L0Memory_43 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  L0Memory_44 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  L0Memory_45 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  L0Memory_46 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  L0Memory_47 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  L0Memory_48 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  L0Memory_49 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  L0Memory_50 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  L0Memory_51 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  L0Memory_52 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  L0Memory_53 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  L0Memory_54 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  L0Memory_55 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  L0Memory_56 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  L0Memory_57 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  L0Memory_58 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  L0Memory_59 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  L0Memory_60 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  L0Memory_61 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  L0Memory_62 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  L0Memory_63 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  L0Memory_64 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  L0Memory_65 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  L0Memory_66 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  L0Memory_67 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  L0Memory_68 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  L0Memory_69 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  L0Memory_70 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  L0Memory_71 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  L0Memory_72 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  L0Memory_73 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  L0Memory_74 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  L0Memory_75 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  L0Memory_76 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  L0Memory_77 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  L0Memory_78 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  L0Memory_79 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  L0Memory_80 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  L0Memory_81 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  L0Memory_82 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  L0Memory_83 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  L0Memory_84 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  L0Memory_85 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  L0Memory_86 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  L0Memory_87 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  L0Memory_88 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  L0Memory_89 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  L0Memory_90 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  L0Memory_91 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  L0Memory_92 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  L0Memory_93 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  L0Memory_94 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  L0Memory_95 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  L0Memory_96 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  L0Memory_97 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  L0Memory_98 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  L0Memory_99 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  state = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  mux2out_reg = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  mux3out_reg = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  count = _RAND_104[9:0];
  _RAND_105 = {1{`RANDOM}};
  count_max = _RAND_105[9:0];
  _RAND_106 = {1{`RANDOM}};
  L0index_begin = _RAND_106[5:0];
  _RAND_107 = {1{`RANDOM}};
  GRU_out_width = _RAND_107[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PE_3(
  input         clock,
  input         reset,
  input  [15:0] io_FromAbovePE,
  input  [15:0] io_FromLeftPE,
  input  [15:0] io_FromL1,
  input  [11:0] io_control_signal_mask,
  output [15:0] io_ToRightPE,
  output [15:0] io_ToBelowPE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] FP16MAC_io_a; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_b; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_c; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_out; // @[PEArray.scala 72:23]
  reg [5:0] L0Index; // @[PEArray.scala 39:24]
  reg [15:0] L0Memory_0; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_1; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_2; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_3; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_4; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_5; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_6; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_7; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_8; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_9; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_10; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_11; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_12; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_13; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_14; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_15; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_16; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_17; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_18; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_19; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_20; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_21; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_22; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_23; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_24; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_25; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_26; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_27; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_28; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_29; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_30; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_31; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_32; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_33; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_34; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_35; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_36; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_37; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_38; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_39; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_40; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_41; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_42; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_43; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_44; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_45; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_46; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_47; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_48; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_49; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_50; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_51; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_52; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_53; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_54; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_55; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_56; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_57; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_58; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_59; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_60; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_61; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_62; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_63; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_64; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_65; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_66; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_67; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_68; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_69; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_70; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_71; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_72; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_73; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_74; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_75; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_76; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_77; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_78; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_79; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_80; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_81; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_82; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_83; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_84; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_85; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_86; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_87; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_88; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_89; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_90; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_91; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_92; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_93; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_94; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_95; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_96; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_97; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_98; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_99; // @[PEArray.scala 40:21]
  reg [2:0] state; // @[PEArray.scala 100:22]
  wire  _T_3 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_12 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_16 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_22 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_31 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_41 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_342 = _T_41 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 231:12 PEArray.scala 32:8]
  wire  _GEN_349 = _T_31 ? 1'h0 : _GEN_342; // @[Conditional.scala 39:67 PEArray.scala 208:12]
  wire  _GEN_459 = _T_22 | _GEN_349; // @[Conditional.scala 39:67 PEArray.scala 32:8]
  wire  _GEN_463 = _T_16 ? 1'h0 : _GEN_459; // @[Conditional.scala 39:67]
  wire  _GEN_572 = _T_12 | _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 149:12]
  wire  sel1 = _T_3 | _GEN_572; // @[Conditional.scala 40:58 PEArray.scala 108:12]
  wire [15:0] MAC_out = FP16MAC_io_out; // @[PEArray.scala 47:21 PEArray.scala 85:11]
  wire  _GEN_465 = _T_16 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 177:12]
  wire  _GEN_580 = _T_12 | _GEN_465; // @[Conditional.scala 39:67 PEArray.scala 34:8]
  wire  sel3 = _T_3 | _GEN_580; // @[Conditional.scala 40:58 PEArray.scala 110:12]
  wire [1:0] _GEN_344 = _T_41 ? 2'h2 : 2'h0; // @[Conditional.scala 39:67 PEArray.scala 233:12 PEArray.scala 35:8]
  wire [1:0] _GEN_351 = _T_31 ? 2'h2 : _GEN_344; // @[Conditional.scala 39:67 PEArray.scala 210:12]
  wire [1:0] _GEN_461 = _T_22 ? 2'h0 : _GEN_351; // @[Conditional.scala 39:67 PEArray.scala 35:8]
  wire [1:0] _GEN_466 = _T_16 ? 2'h0 : _GEN_461; // @[Conditional.scala 39:67 PEArray.scala 178:12]
  wire [1:0] _GEN_574 = _T_12 ? 2'h0 : _GEN_466; // @[Conditional.scala 39:67]
  wire [1:0] sel4 = _T_3 ? 2'h0 : _GEN_574; // @[Conditional.scala 40:58 PEArray.scala 111:12]
  wire [15:0] _GEN_3 = sel4 == 2'h2 ? io_FromL1 : 16'h0; // @[PEArray.scala 65:28 PEArray.scala 66:15 PEArray.scala 69:15]
  wire [15:0] _GEN_4 = sel4 == 2'h1 ? io_FromAbovePE : _GEN_3; // @[PEArray.scala 62:28 PEArray.scala 63:15]
  wire [15:0] mux4out = sel4 == 2'h0 ? 16'h0 : _GEN_4; // @[PEArray.scala 59:22 PEArray.scala 60:13]
  wire [15:0] _GEN_7 = 6'h1 == L0Index ? L0Memory_1 : L0Memory_0; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_8 = 6'h2 == L0Index ? L0Memory_2 : _GEN_7; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_9 = 6'h3 == L0Index ? L0Memory_3 : _GEN_8; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_10 = 6'h4 == L0Index ? L0Memory_4 : _GEN_9; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_11 = 6'h5 == L0Index ? L0Memory_5 : _GEN_10; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_12 = 6'h6 == L0Index ? L0Memory_6 : _GEN_11; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_13 = 6'h7 == L0Index ? L0Memory_7 : _GEN_12; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_14 = 6'h8 == L0Index ? L0Memory_8 : _GEN_13; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_15 = 6'h9 == L0Index ? L0Memory_9 : _GEN_14; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_16 = 6'ha == L0Index ? L0Memory_10 : _GEN_15; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_17 = 6'hb == L0Index ? L0Memory_11 : _GEN_16; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_18 = 6'hc == L0Index ? L0Memory_12 : _GEN_17; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_19 = 6'hd == L0Index ? L0Memory_13 : _GEN_18; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_20 = 6'he == L0Index ? L0Memory_14 : _GEN_19; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_21 = 6'hf == L0Index ? L0Memory_15 : _GEN_20; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_22 = 6'h10 == L0Index ? L0Memory_16 : _GEN_21; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_23 = 6'h11 == L0Index ? L0Memory_17 : _GEN_22; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_24 = 6'h12 == L0Index ? L0Memory_18 : _GEN_23; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_25 = 6'h13 == L0Index ? L0Memory_19 : _GEN_24; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_26 = 6'h14 == L0Index ? L0Memory_20 : _GEN_25; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_27 = 6'h15 == L0Index ? L0Memory_21 : _GEN_26; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_28 = 6'h16 == L0Index ? L0Memory_22 : _GEN_27; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_29 = 6'h17 == L0Index ? L0Memory_23 : _GEN_28; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_30 = 6'h18 == L0Index ? L0Memory_24 : _GEN_29; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_31 = 6'h19 == L0Index ? L0Memory_25 : _GEN_30; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_32 = 6'h1a == L0Index ? L0Memory_26 : _GEN_31; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_33 = 6'h1b == L0Index ? L0Memory_27 : _GEN_32; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_34 = 6'h1c == L0Index ? L0Memory_28 : _GEN_33; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_35 = 6'h1d == L0Index ? L0Memory_29 : _GEN_34; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_36 = 6'h1e == L0Index ? L0Memory_30 : _GEN_35; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_37 = 6'h1f == L0Index ? L0Memory_31 : _GEN_36; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_38 = 6'h20 == L0Index ? L0Memory_32 : _GEN_37; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_39 = 6'h21 == L0Index ? L0Memory_33 : _GEN_38; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_40 = 6'h22 == L0Index ? L0Memory_34 : _GEN_39; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_41 = 6'h23 == L0Index ? L0Memory_35 : _GEN_40; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_42 = 6'h24 == L0Index ? L0Memory_36 : _GEN_41; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_43 = 6'h25 == L0Index ? L0Memory_37 : _GEN_42; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_44 = 6'h26 == L0Index ? L0Memory_38 : _GEN_43; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_45 = 6'h27 == L0Index ? L0Memory_39 : _GEN_44; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_46 = 6'h28 == L0Index ? L0Memory_40 : _GEN_45; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_47 = 6'h29 == L0Index ? L0Memory_41 : _GEN_46; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_48 = 6'h2a == L0Index ? L0Memory_42 : _GEN_47; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_49 = 6'h2b == L0Index ? L0Memory_43 : _GEN_48; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_50 = 6'h2c == L0Index ? L0Memory_44 : _GEN_49; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_51 = 6'h2d == L0Index ? L0Memory_45 : _GEN_50; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_52 = 6'h2e == L0Index ? L0Memory_46 : _GEN_51; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_53 = 6'h2f == L0Index ? L0Memory_47 : _GEN_52; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_54 = 6'h30 == L0Index ? L0Memory_48 : _GEN_53; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_55 = 6'h31 == L0Index ? L0Memory_49 : _GEN_54; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_56 = 6'h32 == L0Index ? L0Memory_50 : _GEN_55; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_57 = 6'h33 == L0Index ? L0Memory_51 : _GEN_56; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_58 = 6'h34 == L0Index ? L0Memory_52 : _GEN_57; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_59 = 6'h35 == L0Index ? L0Memory_53 : _GEN_58; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_60 = 6'h36 == L0Index ? L0Memory_54 : _GEN_59; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_61 = 6'h37 == L0Index ? L0Memory_55 : _GEN_60; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_62 = 6'h38 == L0Index ? L0Memory_56 : _GEN_61; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_63 = 6'h39 == L0Index ? L0Memory_57 : _GEN_62; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_64 = 6'h3a == L0Index ? L0Memory_58 : _GEN_63; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_65 = 6'h3b == L0Index ? L0Memory_59 : _GEN_64; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_66 = 6'h3c == L0Index ? L0Memory_60 : _GEN_65; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_67 = 6'h3d == L0Index ? L0Memory_61 : _GEN_66; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_68 = 6'h3e == L0Index ? L0Memory_62 : _GEN_67; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_69 = 6'h3f == L0Index ? L0Memory_63 : _GEN_68; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [6:0] _GEN_793 = {{1'd0}, L0Index}; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_70 = 7'h40 == _GEN_793 ? L0Memory_64 : _GEN_69; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_71 = 7'h41 == _GEN_793 ? L0Memory_65 : _GEN_70; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_72 = 7'h42 == _GEN_793 ? L0Memory_66 : _GEN_71; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_73 = 7'h43 == _GEN_793 ? L0Memory_67 : _GEN_72; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_74 = 7'h44 == _GEN_793 ? L0Memory_68 : _GEN_73; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_75 = 7'h45 == _GEN_793 ? L0Memory_69 : _GEN_74; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_76 = 7'h46 == _GEN_793 ? L0Memory_70 : _GEN_75; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_77 = 7'h47 == _GEN_793 ? L0Memory_71 : _GEN_76; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_78 = 7'h48 == _GEN_793 ? L0Memory_72 : _GEN_77; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_79 = 7'h49 == _GEN_793 ? L0Memory_73 : _GEN_78; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_80 = 7'h4a == _GEN_793 ? L0Memory_74 : _GEN_79; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_81 = 7'h4b == _GEN_793 ? L0Memory_75 : _GEN_80; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_82 = 7'h4c == _GEN_793 ? L0Memory_76 : _GEN_81; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_83 = 7'h4d == _GEN_793 ? L0Memory_77 : _GEN_82; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_84 = 7'h4e == _GEN_793 ? L0Memory_78 : _GEN_83; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_85 = 7'h4f == _GEN_793 ? L0Memory_79 : _GEN_84; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_86 = 7'h50 == _GEN_793 ? L0Memory_80 : _GEN_85; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_87 = 7'h51 == _GEN_793 ? L0Memory_81 : _GEN_86; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_88 = 7'h52 == _GEN_793 ? L0Memory_82 : _GEN_87; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_89 = 7'h53 == _GEN_793 ? L0Memory_83 : _GEN_88; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_90 = 7'h54 == _GEN_793 ? L0Memory_84 : _GEN_89; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_91 = 7'h55 == _GEN_793 ? L0Memory_85 : _GEN_90; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_92 = 7'h56 == _GEN_793 ? L0Memory_86 : _GEN_91; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_93 = 7'h57 == _GEN_793 ? L0Memory_87 : _GEN_92; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_94 = 7'h58 == _GEN_793 ? L0Memory_88 : _GEN_93; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_95 = 7'h59 == _GEN_793 ? L0Memory_89 : _GEN_94; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_96 = 7'h5a == _GEN_793 ? L0Memory_90 : _GEN_95; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_97 = 7'h5b == _GEN_793 ? L0Memory_91 : _GEN_96; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_98 = 7'h5c == _GEN_793 ? L0Memory_92 : _GEN_97; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_99 = 7'h5d == _GEN_793 ? L0Memory_93 : _GEN_98; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_100 = 7'h5e == _GEN_793 ? L0Memory_94 : _GEN_99; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_101 = 7'h5f == _GEN_793 ? L0Memory_95 : _GEN_100; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_102 = 7'h60 == _GEN_793 ? L0Memory_96 : _GEN_101; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_103 = 7'h61 == _GEN_793 ? L0Memory_97 : _GEN_102; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_104 = 7'h62 == _GEN_793 ? L0Memory_98 : _GEN_103; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_105 = 7'h63 == _GEN_793 ? L0Memory_99 : _GEN_104; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire  _GEN_575 = _T_12 ? 1'h0 : _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 157:12]
  wire  sel5 = _T_3 ? 1'h0 : _GEN_575; // @[Conditional.scala 40:58 PEArray.scala 112:12]
  reg [15:0] mux2out_reg; // @[PEArray.scala 90:28]
  reg [15:0] mux3out_reg; // @[PEArray.scala 91:28]
  reg [9:0] count; // @[PEArray.scala 101:22]
  reg [5:0] GRU_out_width; // @[PEArray.scala 104:26]
  wire [7:0] _GEN_118 = io_control_signal_mask[10] ? 8'h0 : {{2'd0}, GRU_out_width}; // @[PEArray.scala 116:57 PEArray.scala 145:23 PEArray.scala 104:26]
  wire [9:0] _count_T_1 = count + 10'h1; // @[PEArray.scala 162:24]
  wire [9:0] _GEN_120 = count != 10'h33 ? _count_T_1 : count; // @[PEArray.scala 161:27 PEArray.scala 162:15 PEArray.scala 101:22]
  wire [9:0] _GEN_124 = count != 10'h188 ? _count_T_1 : count; // @[PEArray.scala 183:28 PEArray.scala 184:15 PEArray.scala 101:22]
  wire [9:0] _GEN_125 = count == 10'h188 ? 10'h0 : _GEN_124; // @[PEArray.scala 186:28 PEArray.scala 187:15]
  wire [2:0] _GEN_126 = count == 10'h188 ? 3'h0 : state; // @[PEArray.scala 186:28 PEArray.scala 188:15 PEArray.scala 100:22]
  wire [9:0] _GEN_127 = count != 10'h0 ? _count_T_1 : count; // @[PEArray.scala 192:32 PEArray.scala 193:15 PEArray.scala 101:22]
  wire  _T_24 = count == 10'h0; // @[PEArray.scala 195:18]
  wire [5:0] _GEN_128 = count == 10'h0 ? 6'h0 : L0Index; // @[PEArray.scala 195:26 PEArray.scala 196:17 PEArray.scala 39:24]
  wire [9:0] _T_27 = 10'h0 - 10'h1; // @[PEArray.scala 198:51]
  wire [15:0] _GEN_129 = 6'h0 == L0Index ? io_FromL1 : L0Memory_0; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_130 = 6'h1 == L0Index ? io_FromL1 : L0Memory_1; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_131 = 6'h2 == L0Index ? io_FromL1 : L0Memory_2; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_132 = 6'h3 == L0Index ? io_FromL1 : L0Memory_3; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_133 = 6'h4 == L0Index ? io_FromL1 : L0Memory_4; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_134 = 6'h5 == L0Index ? io_FromL1 : L0Memory_5; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_135 = 6'h6 == L0Index ? io_FromL1 : L0Memory_6; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_136 = 6'h7 == L0Index ? io_FromL1 : L0Memory_7; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_137 = 6'h8 == L0Index ? io_FromL1 : L0Memory_8; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_138 = 6'h9 == L0Index ? io_FromL1 : L0Memory_9; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_139 = 6'ha == L0Index ? io_FromL1 : L0Memory_10; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_140 = 6'hb == L0Index ? io_FromL1 : L0Memory_11; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_141 = 6'hc == L0Index ? io_FromL1 : L0Memory_12; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_142 = 6'hd == L0Index ? io_FromL1 : L0Memory_13; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_143 = 6'he == L0Index ? io_FromL1 : L0Memory_14; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_144 = 6'hf == L0Index ? io_FromL1 : L0Memory_15; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_145 = 6'h10 == L0Index ? io_FromL1 : L0Memory_16; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_146 = 6'h11 == L0Index ? io_FromL1 : L0Memory_17; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_147 = 6'h12 == L0Index ? io_FromL1 : L0Memory_18; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_148 = 6'h13 == L0Index ? io_FromL1 : L0Memory_19; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_149 = 6'h14 == L0Index ? io_FromL1 : L0Memory_20; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_150 = 6'h15 == L0Index ? io_FromL1 : L0Memory_21; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_151 = 6'h16 == L0Index ? io_FromL1 : L0Memory_22; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_152 = 6'h17 == L0Index ? io_FromL1 : L0Memory_23; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_153 = 6'h18 == L0Index ? io_FromL1 : L0Memory_24; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_154 = 6'h19 == L0Index ? io_FromL1 : L0Memory_25; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_155 = 6'h1a == L0Index ? io_FromL1 : L0Memory_26; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_156 = 6'h1b == L0Index ? io_FromL1 : L0Memory_27; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_157 = 6'h1c == L0Index ? io_FromL1 : L0Memory_28; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_158 = 6'h1d == L0Index ? io_FromL1 : L0Memory_29; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_159 = 6'h1e == L0Index ? io_FromL1 : L0Memory_30; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_160 = 6'h1f == L0Index ? io_FromL1 : L0Memory_31; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_161 = 6'h20 == L0Index ? io_FromL1 : L0Memory_32; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_162 = 6'h21 == L0Index ? io_FromL1 : L0Memory_33; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_163 = 6'h22 == L0Index ? io_FromL1 : L0Memory_34; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_164 = 6'h23 == L0Index ? io_FromL1 : L0Memory_35; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_165 = 6'h24 == L0Index ? io_FromL1 : L0Memory_36; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_166 = 6'h25 == L0Index ? io_FromL1 : L0Memory_37; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_167 = 6'h26 == L0Index ? io_FromL1 : L0Memory_38; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_168 = 6'h27 == L0Index ? io_FromL1 : L0Memory_39; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_169 = 6'h28 == L0Index ? io_FromL1 : L0Memory_40; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_170 = 6'h29 == L0Index ? io_FromL1 : L0Memory_41; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_171 = 6'h2a == L0Index ? io_FromL1 : L0Memory_42; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_172 = 6'h2b == L0Index ? io_FromL1 : L0Memory_43; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_173 = 6'h2c == L0Index ? io_FromL1 : L0Memory_44; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_174 = 6'h2d == L0Index ? io_FromL1 : L0Memory_45; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_175 = 6'h2e == L0Index ? io_FromL1 : L0Memory_46; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_176 = 6'h2f == L0Index ? io_FromL1 : L0Memory_47; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_177 = 6'h30 == L0Index ? io_FromL1 : L0Memory_48; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_178 = 6'h31 == L0Index ? io_FromL1 : L0Memory_49; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_179 = 6'h32 == L0Index ? io_FromL1 : L0Memory_50; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_180 = 6'h33 == L0Index ? io_FromL1 : L0Memory_51; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_181 = 6'h34 == L0Index ? io_FromL1 : L0Memory_52; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_182 = 6'h35 == L0Index ? io_FromL1 : L0Memory_53; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_183 = 6'h36 == L0Index ? io_FromL1 : L0Memory_54; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_184 = 6'h37 == L0Index ? io_FromL1 : L0Memory_55; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_185 = 6'h38 == L0Index ? io_FromL1 : L0Memory_56; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_186 = 6'h39 == L0Index ? io_FromL1 : L0Memory_57; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_187 = 6'h3a == L0Index ? io_FromL1 : L0Memory_58; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_188 = 6'h3b == L0Index ? io_FromL1 : L0Memory_59; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_189 = 6'h3c == L0Index ? io_FromL1 : L0Memory_60; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_190 = 6'h3d == L0Index ? io_FromL1 : L0Memory_61; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_191 = 6'h3e == L0Index ? io_FromL1 : L0Memory_62; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_192 = 6'h3f == L0Index ? io_FromL1 : L0Memory_63; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_193 = 7'h40 == _GEN_793 ? io_FromL1 : L0Memory_64; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_194 = 7'h41 == _GEN_793 ? io_FromL1 : L0Memory_65; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_195 = 7'h42 == _GEN_793 ? io_FromL1 : L0Memory_66; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_196 = 7'h43 == _GEN_793 ? io_FromL1 : L0Memory_67; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_197 = 7'h44 == _GEN_793 ? io_FromL1 : L0Memory_68; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_198 = 7'h45 == _GEN_793 ? io_FromL1 : L0Memory_69; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_199 = 7'h46 == _GEN_793 ? io_FromL1 : L0Memory_70; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_200 = 7'h47 == _GEN_793 ? io_FromL1 : L0Memory_71; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_201 = 7'h48 == _GEN_793 ? io_FromL1 : L0Memory_72; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_202 = 7'h49 == _GEN_793 ? io_FromL1 : L0Memory_73; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_203 = 7'h4a == _GEN_793 ? io_FromL1 : L0Memory_74; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_204 = 7'h4b == _GEN_793 ? io_FromL1 : L0Memory_75; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_205 = 7'h4c == _GEN_793 ? io_FromL1 : L0Memory_76; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_206 = 7'h4d == _GEN_793 ? io_FromL1 : L0Memory_77; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_207 = 7'h4e == _GEN_793 ? io_FromL1 : L0Memory_78; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_208 = 7'h4f == _GEN_793 ? io_FromL1 : L0Memory_79; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_209 = 7'h50 == _GEN_793 ? io_FromL1 : L0Memory_80; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_210 = 7'h51 == _GEN_793 ? io_FromL1 : L0Memory_81; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_211 = 7'h52 == _GEN_793 ? io_FromL1 : L0Memory_82; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_212 = 7'h53 == _GEN_793 ? io_FromL1 : L0Memory_83; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_213 = 7'h54 == _GEN_793 ? io_FromL1 : L0Memory_84; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_214 = 7'h55 == _GEN_793 ? io_FromL1 : L0Memory_85; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_215 = 7'h56 == _GEN_793 ? io_FromL1 : L0Memory_86; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_216 = 7'h57 == _GEN_793 ? io_FromL1 : L0Memory_87; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_217 = 7'h58 == _GEN_793 ? io_FromL1 : L0Memory_88; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_218 = 7'h59 == _GEN_793 ? io_FromL1 : L0Memory_89; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_219 = 7'h5a == _GEN_793 ? io_FromL1 : L0Memory_90; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_220 = 7'h5b == _GEN_793 ? io_FromL1 : L0Memory_91; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_221 = 7'h5c == _GEN_793 ? io_FromL1 : L0Memory_92; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_222 = 7'h5d == _GEN_793 ? io_FromL1 : L0Memory_93; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_223 = 7'h5e == _GEN_793 ? io_FromL1 : L0Memory_94; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_224 = 7'h5f == _GEN_793 ? io_FromL1 : L0Memory_95; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_225 = 7'h60 == _GEN_793 ? io_FromL1 : L0Memory_96; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_226 = 7'h61 == _GEN_793 ? io_FromL1 : L0Memory_97; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_227 = 7'h62 == _GEN_793 ? io_FromL1 : L0Memory_98; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_228 = 7'h63 == _GEN_793 ? io_FromL1 : L0Memory_99; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [5:0] _L0Index_T_2 = L0Index + 6'h1; // @[PEArray.scala 200:28]
  wire [15:0] _GEN_229 = count >= 10'h1 & count <= _T_27 ? _GEN_129 : L0Memory_0; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_230 = count >= 10'h1 & count <= _T_27 ? _GEN_130 : L0Memory_1; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_231 = count >= 10'h1 & count <= _T_27 ? _GEN_131 : L0Memory_2; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_232 = count >= 10'h1 & count <= _T_27 ? _GEN_132 : L0Memory_3; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_233 = count >= 10'h1 & count <= _T_27 ? _GEN_133 : L0Memory_4; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_234 = count >= 10'h1 & count <= _T_27 ? _GEN_134 : L0Memory_5; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_235 = count >= 10'h1 & count <= _T_27 ? _GEN_135 : L0Memory_6; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_236 = count >= 10'h1 & count <= _T_27 ? _GEN_136 : L0Memory_7; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_237 = count >= 10'h1 & count <= _T_27 ? _GEN_137 : L0Memory_8; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_238 = count >= 10'h1 & count <= _T_27 ? _GEN_138 : L0Memory_9; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_239 = count >= 10'h1 & count <= _T_27 ? _GEN_139 : L0Memory_10; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_240 = count >= 10'h1 & count <= _T_27 ? _GEN_140 : L0Memory_11; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_241 = count >= 10'h1 & count <= _T_27 ? _GEN_141 : L0Memory_12; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_242 = count >= 10'h1 & count <= _T_27 ? _GEN_142 : L0Memory_13; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_243 = count >= 10'h1 & count <= _T_27 ? _GEN_143 : L0Memory_14; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_244 = count >= 10'h1 & count <= _T_27 ? _GEN_144 : L0Memory_15; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_245 = count >= 10'h1 & count <= _T_27 ? _GEN_145 : L0Memory_16; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_246 = count >= 10'h1 & count <= _T_27 ? _GEN_146 : L0Memory_17; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_247 = count >= 10'h1 & count <= _T_27 ? _GEN_147 : L0Memory_18; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_248 = count >= 10'h1 & count <= _T_27 ? _GEN_148 : L0Memory_19; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_249 = count >= 10'h1 & count <= _T_27 ? _GEN_149 : L0Memory_20; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_250 = count >= 10'h1 & count <= _T_27 ? _GEN_150 : L0Memory_21; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_251 = count >= 10'h1 & count <= _T_27 ? _GEN_151 : L0Memory_22; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_252 = count >= 10'h1 & count <= _T_27 ? _GEN_152 : L0Memory_23; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_253 = count >= 10'h1 & count <= _T_27 ? _GEN_153 : L0Memory_24; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_254 = count >= 10'h1 & count <= _T_27 ? _GEN_154 : L0Memory_25; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_255 = count >= 10'h1 & count <= _T_27 ? _GEN_155 : L0Memory_26; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_256 = count >= 10'h1 & count <= _T_27 ? _GEN_156 : L0Memory_27; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_257 = count >= 10'h1 & count <= _T_27 ? _GEN_157 : L0Memory_28; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_258 = count >= 10'h1 & count <= _T_27 ? _GEN_158 : L0Memory_29; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_259 = count >= 10'h1 & count <= _T_27 ? _GEN_159 : L0Memory_30; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_260 = count >= 10'h1 & count <= _T_27 ? _GEN_160 : L0Memory_31; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_261 = count >= 10'h1 & count <= _T_27 ? _GEN_161 : L0Memory_32; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_262 = count >= 10'h1 & count <= _T_27 ? _GEN_162 : L0Memory_33; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_263 = count >= 10'h1 & count <= _T_27 ? _GEN_163 : L0Memory_34; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_264 = count >= 10'h1 & count <= _T_27 ? _GEN_164 : L0Memory_35; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_265 = count >= 10'h1 & count <= _T_27 ? _GEN_165 : L0Memory_36; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_266 = count >= 10'h1 & count <= _T_27 ? _GEN_166 : L0Memory_37; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_267 = count >= 10'h1 & count <= _T_27 ? _GEN_167 : L0Memory_38; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_268 = count >= 10'h1 & count <= _T_27 ? _GEN_168 : L0Memory_39; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_269 = count >= 10'h1 & count <= _T_27 ? _GEN_169 : L0Memory_40; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_270 = count >= 10'h1 & count <= _T_27 ? _GEN_170 : L0Memory_41; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_271 = count >= 10'h1 & count <= _T_27 ? _GEN_171 : L0Memory_42; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_272 = count >= 10'h1 & count <= _T_27 ? _GEN_172 : L0Memory_43; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_273 = count >= 10'h1 & count <= _T_27 ? _GEN_173 : L0Memory_44; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_274 = count >= 10'h1 & count <= _T_27 ? _GEN_174 : L0Memory_45; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_275 = count >= 10'h1 & count <= _T_27 ? _GEN_175 : L0Memory_46; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_276 = count >= 10'h1 & count <= _T_27 ? _GEN_176 : L0Memory_47; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_277 = count >= 10'h1 & count <= _T_27 ? _GEN_177 : L0Memory_48; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_278 = count >= 10'h1 & count <= _T_27 ? _GEN_178 : L0Memory_49; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_279 = count >= 10'h1 & count <= _T_27 ? _GEN_179 : L0Memory_50; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_280 = count >= 10'h1 & count <= _T_27 ? _GEN_180 : L0Memory_51; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_281 = count >= 10'h1 & count <= _T_27 ? _GEN_181 : L0Memory_52; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_282 = count >= 10'h1 & count <= _T_27 ? _GEN_182 : L0Memory_53; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_283 = count >= 10'h1 & count <= _T_27 ? _GEN_183 : L0Memory_54; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_284 = count >= 10'h1 & count <= _T_27 ? _GEN_184 : L0Memory_55; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_285 = count >= 10'h1 & count <= _T_27 ? _GEN_185 : L0Memory_56; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_286 = count >= 10'h1 & count <= _T_27 ? _GEN_186 : L0Memory_57; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_287 = count >= 10'h1 & count <= _T_27 ? _GEN_187 : L0Memory_58; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_288 = count >= 10'h1 & count <= _T_27 ? _GEN_188 : L0Memory_59; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_289 = count >= 10'h1 & count <= _T_27 ? _GEN_189 : L0Memory_60; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_290 = count >= 10'h1 & count <= _T_27 ? _GEN_190 : L0Memory_61; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_291 = count >= 10'h1 & count <= _T_27 ? _GEN_191 : L0Memory_62; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_292 = count >= 10'h1 & count <= _T_27 ? _GEN_192 : L0Memory_63; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_293 = count >= 10'h1 & count <= _T_27 ? _GEN_193 : L0Memory_64; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_294 = count >= 10'h1 & count <= _T_27 ? _GEN_194 : L0Memory_65; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_295 = count >= 10'h1 & count <= _T_27 ? _GEN_195 : L0Memory_66; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_296 = count >= 10'h1 & count <= _T_27 ? _GEN_196 : L0Memory_67; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_297 = count >= 10'h1 & count <= _T_27 ? _GEN_197 : L0Memory_68; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_298 = count >= 10'h1 & count <= _T_27 ? _GEN_198 : L0Memory_69; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_299 = count >= 10'h1 & count <= _T_27 ? _GEN_199 : L0Memory_70; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_300 = count >= 10'h1 & count <= _T_27 ? _GEN_200 : L0Memory_71; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_301 = count >= 10'h1 & count <= _T_27 ? _GEN_201 : L0Memory_72; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_302 = count >= 10'h1 & count <= _T_27 ? _GEN_202 : L0Memory_73; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_303 = count >= 10'h1 & count <= _T_27 ? _GEN_203 : L0Memory_74; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_304 = count >= 10'h1 & count <= _T_27 ? _GEN_204 : L0Memory_75; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_305 = count >= 10'h1 & count <= _T_27 ? _GEN_205 : L0Memory_76; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_306 = count >= 10'h1 & count <= _T_27 ? _GEN_206 : L0Memory_77; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_307 = count >= 10'h1 & count <= _T_27 ? _GEN_207 : L0Memory_78; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_308 = count >= 10'h1 & count <= _T_27 ? _GEN_208 : L0Memory_79; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_309 = count >= 10'h1 & count <= _T_27 ? _GEN_209 : L0Memory_80; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_310 = count >= 10'h1 & count <= _T_27 ? _GEN_210 : L0Memory_81; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_311 = count >= 10'h1 & count <= _T_27 ? _GEN_211 : L0Memory_82; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_312 = count >= 10'h1 & count <= _T_27 ? _GEN_212 : L0Memory_83; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_313 = count >= 10'h1 & count <= _T_27 ? _GEN_213 : L0Memory_84; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_314 = count >= 10'h1 & count <= _T_27 ? _GEN_214 : L0Memory_85; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_315 = count >= 10'h1 & count <= _T_27 ? _GEN_215 : L0Memory_86; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_316 = count >= 10'h1 & count <= _T_27 ? _GEN_216 : L0Memory_87; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_317 = count >= 10'h1 & count <= _T_27 ? _GEN_217 : L0Memory_88; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_318 = count >= 10'h1 & count <= _T_27 ? _GEN_218 : L0Memory_89; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_319 = count >= 10'h1 & count <= _T_27 ? _GEN_219 : L0Memory_90; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_320 = count >= 10'h1 & count <= _T_27 ? _GEN_220 : L0Memory_91; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_321 = count >= 10'h1 & count <= _T_27 ? _GEN_221 : L0Memory_92; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_322 = count >= 10'h1 & count <= _T_27 ? _GEN_222 : L0Memory_93; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_323 = count >= 10'h1 & count <= _T_27 ? _GEN_223 : L0Memory_94; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_324 = count >= 10'h1 & count <= _T_27 ? _GEN_224 : L0Memory_95; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_325 = count >= 10'h1 & count <= _T_27 ? _GEN_225 : L0Memory_96; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_326 = count >= 10'h1 & count <= _T_27 ? _GEN_226 : L0Memory_97; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_327 = count >= 10'h1 & count <= _T_27 ? _GEN_227 : L0Memory_98; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_328 = count >= 10'h1 & count <= _T_27 ? _GEN_228 : L0Memory_99; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [5:0] _GEN_329 = count >= 10'h1 & count <= _T_27 ? _L0Index_T_2 : _GEN_128; // @[PEArray.scala 198:59 PEArray.scala 200:17]
  wire [9:0] _GEN_330 = _T_24 ? 10'h0 : _GEN_127; // @[PEArray.scala 202:32 PEArray.scala 203:15]
  wire [2:0] _GEN_331 = _T_24 ? 3'h0 : state; // @[PEArray.scala 202:32 PEArray.scala 204:15 PEArray.scala 100:22]
  wire [9:0] _GEN_865 = {{4'd0}, GRU_out_width}; // @[PEArray.scala 220:19]
  wire [9:0] _GEN_0 = count % _GEN_865; // @[PEArray.scala 220:19]
  wire [5:0] _T_36 = _GEN_0[5:0]; // @[PEArray.scala 220:19]
  wire [5:0] _T_38 = GRU_out_width - 6'h1; // @[PEArray.scala 220:55]
  wire [5:0] _GEN_334 = _T_36 == _T_38 ? _L0Index_T_2 : 6'h0; // @[PEArray.scala 220:62 PEArray.scala 221:17 PEArray.scala 214:15]
  wire [5:0] _GEN_346 = _T_41 ? _GEN_334 : L0Index; // @[Conditional.scala 39:67 PEArray.scala 39:24]
  wire [9:0] _GEN_347 = _T_41 ? _GEN_330 : count; // @[Conditional.scala 39:67 PEArray.scala 101:22]
  wire [2:0] _GEN_348 = _T_41 ? _GEN_331 : state; // @[Conditional.scala 39:67 PEArray.scala 100:22]
  wire [5:0] _GEN_353 = _T_31 ? _GEN_334 : _GEN_346; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_354 = _T_31 ? _GEN_330 : _GEN_347; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_355 = _T_31 ? _GEN_331 : _GEN_348; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_356 = _T_22 ? _GEN_330 : _GEN_354; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_357 = _T_22 ? _GEN_329 : _GEN_353; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_458 = _T_22 ? _GEN_331 : _GEN_355; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_690 = _T_3 ? _GEN_118 : {{2'd0}, GRU_out_width}; // @[Conditional.scala 40:58 PEArray.scala 104:26]
  FP16MulAdder FP16MAC ( // @[PEArray.scala 72:23]
    .io_a(FP16MAC_io_a),
    .io_b(FP16MAC_io_b),
    .io_c(FP16MAC_io_c),
    .io_out(FP16MAC_io_out)
  );
  assign io_ToRightPE = mux3out_reg; // @[PEArray.scala 95:16]
  assign io_ToBelowPE = mux2out_reg; // @[PEArray.scala 94:16]
  assign FP16MAC_io_a = sel1 ? io_FromL1 : io_FromLeftPE; // @[PEArray.scala 50:14 PEArray.scala 50:23 PEArray.scala 51:24]
  assign FP16MAC_io_b = sel5 ? mux4out : _GEN_105; // @[PEArray.scala 77:13 PEArray.scala 78:18 PEArray.scala 81:18]
  assign FP16MAC_io_c = sel5 ? _GEN_105 : mux4out; // @[PEArray.scala 77:13 PEArray.scala 79:18 PEArray.scala 82:18]
  always @(posedge clock) begin
    if (reset) begin // @[PEArray.scala 39:24]
      L0Index <= 6'h0; // @[PEArray.scala 39:24]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h0; // @[PEArray.scala 159:15]
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h4; // @[PEArray.scala 181:15]
      end else begin
        L0Index <= _GEN_357;
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_0 <= _GEN_229;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_1 <= _GEN_230;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_2 <= _GEN_231;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_3 <= _GEN_232;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_4 <= _GEN_233;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_5 <= _GEN_234;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_6 <= _GEN_235;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_7 <= _GEN_236;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_8 <= _GEN_237;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_9 <= _GEN_238;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_10 <= _GEN_239;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_11 <= _GEN_240;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_12 <= _GEN_241;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_13 <= _GEN_242;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_14 <= _GEN_243;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_15 <= _GEN_244;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_16 <= _GEN_245;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_17 <= _GEN_246;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_18 <= _GEN_247;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_19 <= _GEN_248;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_20 <= _GEN_249;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_21 <= _GEN_250;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_22 <= _GEN_251;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_23 <= _GEN_252;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_24 <= _GEN_253;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_25 <= _GEN_254;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_26 <= _GEN_255;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_27 <= _GEN_256;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_28 <= _GEN_257;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_29 <= _GEN_258;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_30 <= _GEN_259;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_31 <= _GEN_260;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_32 <= _GEN_261;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_33 <= _GEN_262;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_34 <= _GEN_263;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_35 <= _GEN_264;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_36 <= _GEN_265;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_37 <= _GEN_266;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_38 <= _GEN_267;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_39 <= _GEN_268;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_40 <= _GEN_269;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_41 <= _GEN_270;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_42 <= _GEN_271;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_43 <= _GEN_272;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_44 <= _GEN_273;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_45 <= _GEN_274;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_46 <= _GEN_275;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_47 <= _GEN_276;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_48 <= _GEN_277;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_49 <= _GEN_278;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_50 <= _GEN_279;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_51 <= _GEN_280;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_52 <= _GEN_281;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_53 <= _GEN_282;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_54 <= _GEN_283;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_55 <= _GEN_284;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_56 <= _GEN_285;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_57 <= _GEN_286;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_58 <= _GEN_287;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_59 <= _GEN_288;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_60 <= _GEN_289;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_61 <= _GEN_290;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_62 <= _GEN_291;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_63 <= _GEN_292;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_64 <= _GEN_293;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_65 <= _GEN_294;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_66 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_67 <= _GEN_296;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_68 <= _GEN_297;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_69 <= _GEN_298;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_70 <= _GEN_299;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_71 <= _GEN_300;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_72 <= _GEN_301;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_73 <= _GEN_302;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_74 <= _GEN_303;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_75 <= _GEN_304;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_76 <= _GEN_305;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_77 <= _GEN_306;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_78 <= _GEN_307;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_79 <= _GEN_308;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_80 <= _GEN_309;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_81 <= _GEN_310;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_82 <= _GEN_311;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_83 <= _GEN_312;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_84 <= _GEN_313;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_85 <= _GEN_314;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_86 <= _GEN_315;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_87 <= _GEN_316;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_88 <= _GEN_317;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_89 <= _GEN_318;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_90 <= _GEN_319;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_91 <= _GEN_320;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_92 <= _GEN_321;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_93 <= _GEN_322;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_94 <= _GEN_323;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_95 <= _GEN_324;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_96 <= _GEN_325;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_97 <= _GEN_326;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_98 <= _GEN_327;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_99 <= _GEN_328;
          end
        end
      end
    end
    if (reset) begin // @[PEArray.scala 100:22]
      state <= 3'h0; // @[PEArray.scala 100:22]
    end else if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[10]) begin // @[PEArray.scala 116:57]
        state <= 3'h1;
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      if (count == 10'h33) begin // @[PEArray.scala 164:27]
        state <= 3'h0; // @[PEArray.scala 166:15]
      end
    end else if (_T_16) begin // @[Conditional.scala 39:67]
      state <= _GEN_126;
    end else begin
      state <= _GEN_458;
    end
    if (reset) begin // @[PEArray.scala 90:28]
      mux2out_reg <= 16'h0; // @[PEArray.scala 90:28]
    end else begin
      mux2out_reg <= MAC_out; // @[PEArray.scala 90:28]
    end
    if (reset) begin // @[PEArray.scala 91:28]
      mux3out_reg <= 16'h0; // @[PEArray.scala 91:28]
    end else if (sel3) begin // @[PEArray.scala 56:14]
      mux3out_reg <= MAC_out; // @[PEArray.scala 56:23]
    end else if (sel1) begin // @[PEArray.scala 50:14]
      mux3out_reg <= io_FromL1; // @[PEArray.scala 50:23]
    end else begin
      mux3out_reg <= io_FromLeftPE; // @[PEArray.scala 51:24]
    end
    if (reset) begin // @[PEArray.scala 101:22]
      count <= 10'h0; // @[PEArray.scala 101:22]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        if (count == 10'h33) begin // @[PEArray.scala 164:27]
          count <= 10'h0; // @[PEArray.scala 165:15]
        end else begin
          count <= _GEN_120;
        end
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        count <= _GEN_125;
      end else begin
        count <= _GEN_356;
      end
    end
    GRU_out_width <= _GEN_690[5:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  L0Index = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  L0Memory_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  L0Memory_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  L0Memory_2 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  L0Memory_3 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  L0Memory_4 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  L0Memory_5 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  L0Memory_6 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  L0Memory_7 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  L0Memory_8 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  L0Memory_9 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  L0Memory_10 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  L0Memory_11 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  L0Memory_12 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  L0Memory_13 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  L0Memory_14 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  L0Memory_15 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  L0Memory_16 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  L0Memory_17 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  L0Memory_18 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  L0Memory_19 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  L0Memory_20 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  L0Memory_21 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  L0Memory_22 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  L0Memory_23 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  L0Memory_24 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  L0Memory_25 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  L0Memory_26 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  L0Memory_27 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  L0Memory_28 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  L0Memory_29 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  L0Memory_30 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  L0Memory_31 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  L0Memory_32 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  L0Memory_33 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  L0Memory_34 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  L0Memory_35 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  L0Memory_36 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  L0Memory_37 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  L0Memory_38 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  L0Memory_39 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  L0Memory_40 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  L0Memory_41 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  L0Memory_42 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  L0Memory_43 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  L0Memory_44 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  L0Memory_45 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  L0Memory_46 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  L0Memory_47 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  L0Memory_48 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  L0Memory_49 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  L0Memory_50 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  L0Memory_51 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  L0Memory_52 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  L0Memory_53 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  L0Memory_54 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  L0Memory_55 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  L0Memory_56 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  L0Memory_57 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  L0Memory_58 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  L0Memory_59 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  L0Memory_60 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  L0Memory_61 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  L0Memory_62 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  L0Memory_63 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  L0Memory_64 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  L0Memory_65 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  L0Memory_66 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  L0Memory_67 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  L0Memory_68 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  L0Memory_69 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  L0Memory_70 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  L0Memory_71 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  L0Memory_72 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  L0Memory_73 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  L0Memory_74 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  L0Memory_75 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  L0Memory_76 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  L0Memory_77 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  L0Memory_78 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  L0Memory_79 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  L0Memory_80 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  L0Memory_81 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  L0Memory_82 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  L0Memory_83 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  L0Memory_84 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  L0Memory_85 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  L0Memory_86 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  L0Memory_87 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  L0Memory_88 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  L0Memory_89 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  L0Memory_90 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  L0Memory_91 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  L0Memory_92 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  L0Memory_93 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  L0Memory_94 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  L0Memory_95 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  L0Memory_96 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  L0Memory_97 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  L0Memory_98 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  L0Memory_99 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  state = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  mux2out_reg = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  mux3out_reg = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  count = _RAND_104[9:0];
  _RAND_105 = {1{`RANDOM}};
  GRU_out_width = _RAND_105[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PE_4(
  input         clock,
  input         reset,
  input  [15:0] io_FromAbovePE,
  input  [15:0] io_FromLeftPE,
  input  [15:0] io_FromL1,
  input  [11:0] io_control_signal_mask,
  output [15:0] io_ToRightPE,
  output [15:0] io_ToBelowPE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] FP16MAC_io_a; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_b; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_c; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_out; // @[PEArray.scala 72:23]
  reg [5:0] L0Index; // @[PEArray.scala 39:24]
  reg [15:0] L0Memory_0; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_1; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_2; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_3; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_4; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_5; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_6; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_7; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_8; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_9; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_10; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_11; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_12; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_13; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_14; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_15; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_16; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_17; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_18; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_19; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_20; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_21; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_22; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_23; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_24; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_25; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_26; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_27; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_28; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_29; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_30; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_31; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_32; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_33; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_34; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_35; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_36; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_37; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_38; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_39; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_40; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_41; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_42; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_43; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_44; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_45; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_46; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_47; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_48; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_49; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_50; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_51; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_52; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_53; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_54; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_55; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_56; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_57; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_58; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_59; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_60; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_61; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_62; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_63; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_64; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_65; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_66; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_67; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_68; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_69; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_70; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_71; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_72; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_73; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_74; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_75; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_76; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_77; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_78; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_79; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_80; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_81; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_82; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_83; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_84; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_85; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_86; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_87; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_88; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_89; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_90; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_91; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_92; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_93; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_94; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_95; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_96; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_97; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_98; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_99; // @[PEArray.scala 40:21]
  reg [2:0] state; // @[PEArray.scala 100:22]
  wire  _T_3 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_12 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_16 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_22 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_31 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_41 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_342 = _T_41 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 231:12 PEArray.scala 32:8]
  wire  _GEN_349 = _T_31 ? 1'h0 : _GEN_342; // @[Conditional.scala 39:67 PEArray.scala 208:12]
  wire  _GEN_459 = _T_22 | _GEN_349; // @[Conditional.scala 39:67 PEArray.scala 32:8]
  wire  _GEN_463 = _T_16 ? 1'h0 : _GEN_459; // @[Conditional.scala 39:67]
  wire  _GEN_572 = _T_12 | _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 149:12]
  wire  sel1 = _T_3 | _GEN_572; // @[Conditional.scala 40:58 PEArray.scala 108:12]
  wire [15:0] MAC_out = FP16MAC_io_out; // @[PEArray.scala 47:21 PEArray.scala 85:11]
  wire  _GEN_465 = _T_16 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 177:12]
  wire  _GEN_580 = _T_12 | _GEN_465; // @[Conditional.scala 39:67 PEArray.scala 34:8]
  wire  sel3 = _T_3 | _GEN_580; // @[Conditional.scala 40:58 PEArray.scala 110:12]
  wire [1:0] _GEN_344 = _T_41 ? 2'h2 : 2'h0; // @[Conditional.scala 39:67 PEArray.scala 233:12 PEArray.scala 35:8]
  wire [1:0] _GEN_351 = _T_31 ? 2'h2 : _GEN_344; // @[Conditional.scala 39:67 PEArray.scala 210:12]
  wire [1:0] _GEN_461 = _T_22 ? 2'h0 : _GEN_351; // @[Conditional.scala 39:67 PEArray.scala 35:8]
  wire [1:0] _GEN_466 = _T_16 ? 2'h0 : _GEN_461; // @[Conditional.scala 39:67 PEArray.scala 178:12]
  wire [1:0] _GEN_574 = _T_12 ? 2'h1 : _GEN_466; // @[Conditional.scala 39:67]
  wire [1:0] sel4 = _T_3 ? 2'h0 : _GEN_574; // @[Conditional.scala 40:58 PEArray.scala 111:12]
  wire [15:0] _GEN_3 = sel4 == 2'h2 ? io_FromL1 : 16'h0; // @[PEArray.scala 65:28 PEArray.scala 66:15 PEArray.scala 69:15]
  wire [15:0] _GEN_4 = sel4 == 2'h1 ? io_FromAbovePE : _GEN_3; // @[PEArray.scala 62:28 PEArray.scala 63:15]
  wire [15:0] mux4out = sel4 == 2'h0 ? 16'h0 : _GEN_4; // @[PEArray.scala 59:22 PEArray.scala 60:13]
  wire [15:0] _GEN_7 = 6'h1 == L0Index ? L0Memory_1 : L0Memory_0; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_8 = 6'h2 == L0Index ? L0Memory_2 : _GEN_7; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_9 = 6'h3 == L0Index ? L0Memory_3 : _GEN_8; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_10 = 6'h4 == L0Index ? L0Memory_4 : _GEN_9; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_11 = 6'h5 == L0Index ? L0Memory_5 : _GEN_10; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_12 = 6'h6 == L0Index ? L0Memory_6 : _GEN_11; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_13 = 6'h7 == L0Index ? L0Memory_7 : _GEN_12; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_14 = 6'h8 == L0Index ? L0Memory_8 : _GEN_13; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_15 = 6'h9 == L0Index ? L0Memory_9 : _GEN_14; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_16 = 6'ha == L0Index ? L0Memory_10 : _GEN_15; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_17 = 6'hb == L0Index ? L0Memory_11 : _GEN_16; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_18 = 6'hc == L0Index ? L0Memory_12 : _GEN_17; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_19 = 6'hd == L0Index ? L0Memory_13 : _GEN_18; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_20 = 6'he == L0Index ? L0Memory_14 : _GEN_19; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_21 = 6'hf == L0Index ? L0Memory_15 : _GEN_20; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_22 = 6'h10 == L0Index ? L0Memory_16 : _GEN_21; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_23 = 6'h11 == L0Index ? L0Memory_17 : _GEN_22; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_24 = 6'h12 == L0Index ? L0Memory_18 : _GEN_23; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_25 = 6'h13 == L0Index ? L0Memory_19 : _GEN_24; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_26 = 6'h14 == L0Index ? L0Memory_20 : _GEN_25; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_27 = 6'h15 == L0Index ? L0Memory_21 : _GEN_26; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_28 = 6'h16 == L0Index ? L0Memory_22 : _GEN_27; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_29 = 6'h17 == L0Index ? L0Memory_23 : _GEN_28; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_30 = 6'h18 == L0Index ? L0Memory_24 : _GEN_29; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_31 = 6'h19 == L0Index ? L0Memory_25 : _GEN_30; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_32 = 6'h1a == L0Index ? L0Memory_26 : _GEN_31; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_33 = 6'h1b == L0Index ? L0Memory_27 : _GEN_32; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_34 = 6'h1c == L0Index ? L0Memory_28 : _GEN_33; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_35 = 6'h1d == L0Index ? L0Memory_29 : _GEN_34; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_36 = 6'h1e == L0Index ? L0Memory_30 : _GEN_35; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_37 = 6'h1f == L0Index ? L0Memory_31 : _GEN_36; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_38 = 6'h20 == L0Index ? L0Memory_32 : _GEN_37; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_39 = 6'h21 == L0Index ? L0Memory_33 : _GEN_38; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_40 = 6'h22 == L0Index ? L0Memory_34 : _GEN_39; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_41 = 6'h23 == L0Index ? L0Memory_35 : _GEN_40; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_42 = 6'h24 == L0Index ? L0Memory_36 : _GEN_41; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_43 = 6'h25 == L0Index ? L0Memory_37 : _GEN_42; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_44 = 6'h26 == L0Index ? L0Memory_38 : _GEN_43; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_45 = 6'h27 == L0Index ? L0Memory_39 : _GEN_44; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_46 = 6'h28 == L0Index ? L0Memory_40 : _GEN_45; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_47 = 6'h29 == L0Index ? L0Memory_41 : _GEN_46; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_48 = 6'h2a == L0Index ? L0Memory_42 : _GEN_47; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_49 = 6'h2b == L0Index ? L0Memory_43 : _GEN_48; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_50 = 6'h2c == L0Index ? L0Memory_44 : _GEN_49; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_51 = 6'h2d == L0Index ? L0Memory_45 : _GEN_50; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_52 = 6'h2e == L0Index ? L0Memory_46 : _GEN_51; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_53 = 6'h2f == L0Index ? L0Memory_47 : _GEN_52; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_54 = 6'h30 == L0Index ? L0Memory_48 : _GEN_53; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_55 = 6'h31 == L0Index ? L0Memory_49 : _GEN_54; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_56 = 6'h32 == L0Index ? L0Memory_50 : _GEN_55; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_57 = 6'h33 == L0Index ? L0Memory_51 : _GEN_56; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_58 = 6'h34 == L0Index ? L0Memory_52 : _GEN_57; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_59 = 6'h35 == L0Index ? L0Memory_53 : _GEN_58; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_60 = 6'h36 == L0Index ? L0Memory_54 : _GEN_59; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_61 = 6'h37 == L0Index ? L0Memory_55 : _GEN_60; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_62 = 6'h38 == L0Index ? L0Memory_56 : _GEN_61; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_63 = 6'h39 == L0Index ? L0Memory_57 : _GEN_62; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_64 = 6'h3a == L0Index ? L0Memory_58 : _GEN_63; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_65 = 6'h3b == L0Index ? L0Memory_59 : _GEN_64; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_66 = 6'h3c == L0Index ? L0Memory_60 : _GEN_65; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_67 = 6'h3d == L0Index ? L0Memory_61 : _GEN_66; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_68 = 6'h3e == L0Index ? L0Memory_62 : _GEN_67; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_69 = 6'h3f == L0Index ? L0Memory_63 : _GEN_68; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [6:0] _GEN_793 = {{1'd0}, L0Index}; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_70 = 7'h40 == _GEN_793 ? L0Memory_64 : _GEN_69; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_71 = 7'h41 == _GEN_793 ? L0Memory_65 : _GEN_70; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_72 = 7'h42 == _GEN_793 ? L0Memory_66 : _GEN_71; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_73 = 7'h43 == _GEN_793 ? L0Memory_67 : _GEN_72; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_74 = 7'h44 == _GEN_793 ? L0Memory_68 : _GEN_73; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_75 = 7'h45 == _GEN_793 ? L0Memory_69 : _GEN_74; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_76 = 7'h46 == _GEN_793 ? L0Memory_70 : _GEN_75; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_77 = 7'h47 == _GEN_793 ? L0Memory_71 : _GEN_76; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_78 = 7'h48 == _GEN_793 ? L0Memory_72 : _GEN_77; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_79 = 7'h49 == _GEN_793 ? L0Memory_73 : _GEN_78; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_80 = 7'h4a == _GEN_793 ? L0Memory_74 : _GEN_79; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_81 = 7'h4b == _GEN_793 ? L0Memory_75 : _GEN_80; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_82 = 7'h4c == _GEN_793 ? L0Memory_76 : _GEN_81; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_83 = 7'h4d == _GEN_793 ? L0Memory_77 : _GEN_82; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_84 = 7'h4e == _GEN_793 ? L0Memory_78 : _GEN_83; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_85 = 7'h4f == _GEN_793 ? L0Memory_79 : _GEN_84; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_86 = 7'h50 == _GEN_793 ? L0Memory_80 : _GEN_85; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_87 = 7'h51 == _GEN_793 ? L0Memory_81 : _GEN_86; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_88 = 7'h52 == _GEN_793 ? L0Memory_82 : _GEN_87; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_89 = 7'h53 == _GEN_793 ? L0Memory_83 : _GEN_88; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_90 = 7'h54 == _GEN_793 ? L0Memory_84 : _GEN_89; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_91 = 7'h55 == _GEN_793 ? L0Memory_85 : _GEN_90; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_92 = 7'h56 == _GEN_793 ? L0Memory_86 : _GEN_91; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_93 = 7'h57 == _GEN_793 ? L0Memory_87 : _GEN_92; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_94 = 7'h58 == _GEN_793 ? L0Memory_88 : _GEN_93; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_95 = 7'h59 == _GEN_793 ? L0Memory_89 : _GEN_94; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_96 = 7'h5a == _GEN_793 ? L0Memory_90 : _GEN_95; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_97 = 7'h5b == _GEN_793 ? L0Memory_91 : _GEN_96; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_98 = 7'h5c == _GEN_793 ? L0Memory_92 : _GEN_97; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_99 = 7'h5d == _GEN_793 ? L0Memory_93 : _GEN_98; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_100 = 7'h5e == _GEN_793 ? L0Memory_94 : _GEN_99; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_101 = 7'h5f == _GEN_793 ? L0Memory_95 : _GEN_100; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_102 = 7'h60 == _GEN_793 ? L0Memory_96 : _GEN_101; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_103 = 7'h61 == _GEN_793 ? L0Memory_97 : _GEN_102; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_104 = 7'h62 == _GEN_793 ? L0Memory_98 : _GEN_103; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_105 = 7'h63 == _GEN_793 ? L0Memory_99 : _GEN_104; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire  _GEN_575 = _T_12 ? 1'h0 : _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 157:12]
  wire  sel5 = _T_3 ? 1'h0 : _GEN_575; // @[Conditional.scala 40:58 PEArray.scala 112:12]
  reg [15:0] mux2out_reg; // @[PEArray.scala 90:28]
  reg [15:0] mux3out_reg; // @[PEArray.scala 91:28]
  reg [9:0] count; // @[PEArray.scala 101:22]
  reg [5:0] GRU_out_width; // @[PEArray.scala 104:26]
  wire [7:0] _GEN_118 = io_control_signal_mask[10] ? 8'h0 : {{2'd0}, GRU_out_width}; // @[PEArray.scala 116:57 PEArray.scala 145:23 PEArray.scala 104:26]
  wire [9:0] _count_T_1 = count + 10'h1; // @[PEArray.scala 162:24]
  wire [9:0] _GEN_120 = count != 10'h33 ? _count_T_1 : count; // @[PEArray.scala 161:27 PEArray.scala 162:15 PEArray.scala 101:22]
  wire [9:0] _GEN_124 = count != 10'h188 ? _count_T_1 : count; // @[PEArray.scala 183:28 PEArray.scala 184:15 PEArray.scala 101:22]
  wire [9:0] _GEN_125 = count == 10'h188 ? 10'h0 : _GEN_124; // @[PEArray.scala 186:28 PEArray.scala 187:15]
  wire [2:0] _GEN_126 = count == 10'h188 ? 3'h0 : state; // @[PEArray.scala 186:28 PEArray.scala 188:15 PEArray.scala 100:22]
  wire [9:0] _GEN_127 = count != 10'h0 ? _count_T_1 : count; // @[PEArray.scala 192:32 PEArray.scala 193:15 PEArray.scala 101:22]
  wire  _T_24 = count == 10'h0; // @[PEArray.scala 195:18]
  wire [5:0] _GEN_128 = count == 10'h0 ? 6'h0 : L0Index; // @[PEArray.scala 195:26 PEArray.scala 196:17 PEArray.scala 39:24]
  wire [9:0] _T_27 = 10'h0 - 10'h1; // @[PEArray.scala 198:51]
  wire [15:0] _GEN_129 = 6'h0 == L0Index ? io_FromL1 : L0Memory_0; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_130 = 6'h1 == L0Index ? io_FromL1 : L0Memory_1; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_131 = 6'h2 == L0Index ? io_FromL1 : L0Memory_2; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_132 = 6'h3 == L0Index ? io_FromL1 : L0Memory_3; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_133 = 6'h4 == L0Index ? io_FromL1 : L0Memory_4; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_134 = 6'h5 == L0Index ? io_FromL1 : L0Memory_5; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_135 = 6'h6 == L0Index ? io_FromL1 : L0Memory_6; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_136 = 6'h7 == L0Index ? io_FromL1 : L0Memory_7; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_137 = 6'h8 == L0Index ? io_FromL1 : L0Memory_8; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_138 = 6'h9 == L0Index ? io_FromL1 : L0Memory_9; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_139 = 6'ha == L0Index ? io_FromL1 : L0Memory_10; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_140 = 6'hb == L0Index ? io_FromL1 : L0Memory_11; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_141 = 6'hc == L0Index ? io_FromL1 : L0Memory_12; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_142 = 6'hd == L0Index ? io_FromL1 : L0Memory_13; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_143 = 6'he == L0Index ? io_FromL1 : L0Memory_14; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_144 = 6'hf == L0Index ? io_FromL1 : L0Memory_15; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_145 = 6'h10 == L0Index ? io_FromL1 : L0Memory_16; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_146 = 6'h11 == L0Index ? io_FromL1 : L0Memory_17; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_147 = 6'h12 == L0Index ? io_FromL1 : L0Memory_18; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_148 = 6'h13 == L0Index ? io_FromL1 : L0Memory_19; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_149 = 6'h14 == L0Index ? io_FromL1 : L0Memory_20; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_150 = 6'h15 == L0Index ? io_FromL1 : L0Memory_21; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_151 = 6'h16 == L0Index ? io_FromL1 : L0Memory_22; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_152 = 6'h17 == L0Index ? io_FromL1 : L0Memory_23; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_153 = 6'h18 == L0Index ? io_FromL1 : L0Memory_24; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_154 = 6'h19 == L0Index ? io_FromL1 : L0Memory_25; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_155 = 6'h1a == L0Index ? io_FromL1 : L0Memory_26; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_156 = 6'h1b == L0Index ? io_FromL1 : L0Memory_27; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_157 = 6'h1c == L0Index ? io_FromL1 : L0Memory_28; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_158 = 6'h1d == L0Index ? io_FromL1 : L0Memory_29; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_159 = 6'h1e == L0Index ? io_FromL1 : L0Memory_30; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_160 = 6'h1f == L0Index ? io_FromL1 : L0Memory_31; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_161 = 6'h20 == L0Index ? io_FromL1 : L0Memory_32; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_162 = 6'h21 == L0Index ? io_FromL1 : L0Memory_33; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_163 = 6'h22 == L0Index ? io_FromL1 : L0Memory_34; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_164 = 6'h23 == L0Index ? io_FromL1 : L0Memory_35; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_165 = 6'h24 == L0Index ? io_FromL1 : L0Memory_36; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_166 = 6'h25 == L0Index ? io_FromL1 : L0Memory_37; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_167 = 6'h26 == L0Index ? io_FromL1 : L0Memory_38; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_168 = 6'h27 == L0Index ? io_FromL1 : L0Memory_39; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_169 = 6'h28 == L0Index ? io_FromL1 : L0Memory_40; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_170 = 6'h29 == L0Index ? io_FromL1 : L0Memory_41; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_171 = 6'h2a == L0Index ? io_FromL1 : L0Memory_42; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_172 = 6'h2b == L0Index ? io_FromL1 : L0Memory_43; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_173 = 6'h2c == L0Index ? io_FromL1 : L0Memory_44; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_174 = 6'h2d == L0Index ? io_FromL1 : L0Memory_45; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_175 = 6'h2e == L0Index ? io_FromL1 : L0Memory_46; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_176 = 6'h2f == L0Index ? io_FromL1 : L0Memory_47; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_177 = 6'h30 == L0Index ? io_FromL1 : L0Memory_48; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_178 = 6'h31 == L0Index ? io_FromL1 : L0Memory_49; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_179 = 6'h32 == L0Index ? io_FromL1 : L0Memory_50; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_180 = 6'h33 == L0Index ? io_FromL1 : L0Memory_51; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_181 = 6'h34 == L0Index ? io_FromL1 : L0Memory_52; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_182 = 6'h35 == L0Index ? io_FromL1 : L0Memory_53; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_183 = 6'h36 == L0Index ? io_FromL1 : L0Memory_54; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_184 = 6'h37 == L0Index ? io_FromL1 : L0Memory_55; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_185 = 6'h38 == L0Index ? io_FromL1 : L0Memory_56; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_186 = 6'h39 == L0Index ? io_FromL1 : L0Memory_57; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_187 = 6'h3a == L0Index ? io_FromL1 : L0Memory_58; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_188 = 6'h3b == L0Index ? io_FromL1 : L0Memory_59; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_189 = 6'h3c == L0Index ? io_FromL1 : L0Memory_60; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_190 = 6'h3d == L0Index ? io_FromL1 : L0Memory_61; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_191 = 6'h3e == L0Index ? io_FromL1 : L0Memory_62; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_192 = 6'h3f == L0Index ? io_FromL1 : L0Memory_63; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_193 = 7'h40 == _GEN_793 ? io_FromL1 : L0Memory_64; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_194 = 7'h41 == _GEN_793 ? io_FromL1 : L0Memory_65; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_195 = 7'h42 == _GEN_793 ? io_FromL1 : L0Memory_66; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_196 = 7'h43 == _GEN_793 ? io_FromL1 : L0Memory_67; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_197 = 7'h44 == _GEN_793 ? io_FromL1 : L0Memory_68; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_198 = 7'h45 == _GEN_793 ? io_FromL1 : L0Memory_69; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_199 = 7'h46 == _GEN_793 ? io_FromL1 : L0Memory_70; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_200 = 7'h47 == _GEN_793 ? io_FromL1 : L0Memory_71; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_201 = 7'h48 == _GEN_793 ? io_FromL1 : L0Memory_72; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_202 = 7'h49 == _GEN_793 ? io_FromL1 : L0Memory_73; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_203 = 7'h4a == _GEN_793 ? io_FromL1 : L0Memory_74; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_204 = 7'h4b == _GEN_793 ? io_FromL1 : L0Memory_75; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_205 = 7'h4c == _GEN_793 ? io_FromL1 : L0Memory_76; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_206 = 7'h4d == _GEN_793 ? io_FromL1 : L0Memory_77; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_207 = 7'h4e == _GEN_793 ? io_FromL1 : L0Memory_78; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_208 = 7'h4f == _GEN_793 ? io_FromL1 : L0Memory_79; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_209 = 7'h50 == _GEN_793 ? io_FromL1 : L0Memory_80; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_210 = 7'h51 == _GEN_793 ? io_FromL1 : L0Memory_81; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_211 = 7'h52 == _GEN_793 ? io_FromL1 : L0Memory_82; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_212 = 7'h53 == _GEN_793 ? io_FromL1 : L0Memory_83; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_213 = 7'h54 == _GEN_793 ? io_FromL1 : L0Memory_84; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_214 = 7'h55 == _GEN_793 ? io_FromL1 : L0Memory_85; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_215 = 7'h56 == _GEN_793 ? io_FromL1 : L0Memory_86; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_216 = 7'h57 == _GEN_793 ? io_FromL1 : L0Memory_87; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_217 = 7'h58 == _GEN_793 ? io_FromL1 : L0Memory_88; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_218 = 7'h59 == _GEN_793 ? io_FromL1 : L0Memory_89; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_219 = 7'h5a == _GEN_793 ? io_FromL1 : L0Memory_90; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_220 = 7'h5b == _GEN_793 ? io_FromL1 : L0Memory_91; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_221 = 7'h5c == _GEN_793 ? io_FromL1 : L0Memory_92; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_222 = 7'h5d == _GEN_793 ? io_FromL1 : L0Memory_93; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_223 = 7'h5e == _GEN_793 ? io_FromL1 : L0Memory_94; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_224 = 7'h5f == _GEN_793 ? io_FromL1 : L0Memory_95; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_225 = 7'h60 == _GEN_793 ? io_FromL1 : L0Memory_96; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_226 = 7'h61 == _GEN_793 ? io_FromL1 : L0Memory_97; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_227 = 7'h62 == _GEN_793 ? io_FromL1 : L0Memory_98; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_228 = 7'h63 == _GEN_793 ? io_FromL1 : L0Memory_99; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [5:0] _L0Index_T_2 = L0Index + 6'h1; // @[PEArray.scala 200:28]
  wire [15:0] _GEN_229 = count >= 10'h1 & count <= _T_27 ? _GEN_129 : L0Memory_0; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_230 = count >= 10'h1 & count <= _T_27 ? _GEN_130 : L0Memory_1; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_231 = count >= 10'h1 & count <= _T_27 ? _GEN_131 : L0Memory_2; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_232 = count >= 10'h1 & count <= _T_27 ? _GEN_132 : L0Memory_3; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_233 = count >= 10'h1 & count <= _T_27 ? _GEN_133 : L0Memory_4; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_234 = count >= 10'h1 & count <= _T_27 ? _GEN_134 : L0Memory_5; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_235 = count >= 10'h1 & count <= _T_27 ? _GEN_135 : L0Memory_6; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_236 = count >= 10'h1 & count <= _T_27 ? _GEN_136 : L0Memory_7; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_237 = count >= 10'h1 & count <= _T_27 ? _GEN_137 : L0Memory_8; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_238 = count >= 10'h1 & count <= _T_27 ? _GEN_138 : L0Memory_9; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_239 = count >= 10'h1 & count <= _T_27 ? _GEN_139 : L0Memory_10; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_240 = count >= 10'h1 & count <= _T_27 ? _GEN_140 : L0Memory_11; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_241 = count >= 10'h1 & count <= _T_27 ? _GEN_141 : L0Memory_12; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_242 = count >= 10'h1 & count <= _T_27 ? _GEN_142 : L0Memory_13; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_243 = count >= 10'h1 & count <= _T_27 ? _GEN_143 : L0Memory_14; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_244 = count >= 10'h1 & count <= _T_27 ? _GEN_144 : L0Memory_15; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_245 = count >= 10'h1 & count <= _T_27 ? _GEN_145 : L0Memory_16; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_246 = count >= 10'h1 & count <= _T_27 ? _GEN_146 : L0Memory_17; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_247 = count >= 10'h1 & count <= _T_27 ? _GEN_147 : L0Memory_18; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_248 = count >= 10'h1 & count <= _T_27 ? _GEN_148 : L0Memory_19; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_249 = count >= 10'h1 & count <= _T_27 ? _GEN_149 : L0Memory_20; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_250 = count >= 10'h1 & count <= _T_27 ? _GEN_150 : L0Memory_21; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_251 = count >= 10'h1 & count <= _T_27 ? _GEN_151 : L0Memory_22; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_252 = count >= 10'h1 & count <= _T_27 ? _GEN_152 : L0Memory_23; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_253 = count >= 10'h1 & count <= _T_27 ? _GEN_153 : L0Memory_24; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_254 = count >= 10'h1 & count <= _T_27 ? _GEN_154 : L0Memory_25; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_255 = count >= 10'h1 & count <= _T_27 ? _GEN_155 : L0Memory_26; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_256 = count >= 10'h1 & count <= _T_27 ? _GEN_156 : L0Memory_27; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_257 = count >= 10'h1 & count <= _T_27 ? _GEN_157 : L0Memory_28; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_258 = count >= 10'h1 & count <= _T_27 ? _GEN_158 : L0Memory_29; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_259 = count >= 10'h1 & count <= _T_27 ? _GEN_159 : L0Memory_30; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_260 = count >= 10'h1 & count <= _T_27 ? _GEN_160 : L0Memory_31; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_261 = count >= 10'h1 & count <= _T_27 ? _GEN_161 : L0Memory_32; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_262 = count >= 10'h1 & count <= _T_27 ? _GEN_162 : L0Memory_33; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_263 = count >= 10'h1 & count <= _T_27 ? _GEN_163 : L0Memory_34; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_264 = count >= 10'h1 & count <= _T_27 ? _GEN_164 : L0Memory_35; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_265 = count >= 10'h1 & count <= _T_27 ? _GEN_165 : L0Memory_36; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_266 = count >= 10'h1 & count <= _T_27 ? _GEN_166 : L0Memory_37; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_267 = count >= 10'h1 & count <= _T_27 ? _GEN_167 : L0Memory_38; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_268 = count >= 10'h1 & count <= _T_27 ? _GEN_168 : L0Memory_39; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_269 = count >= 10'h1 & count <= _T_27 ? _GEN_169 : L0Memory_40; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_270 = count >= 10'h1 & count <= _T_27 ? _GEN_170 : L0Memory_41; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_271 = count >= 10'h1 & count <= _T_27 ? _GEN_171 : L0Memory_42; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_272 = count >= 10'h1 & count <= _T_27 ? _GEN_172 : L0Memory_43; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_273 = count >= 10'h1 & count <= _T_27 ? _GEN_173 : L0Memory_44; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_274 = count >= 10'h1 & count <= _T_27 ? _GEN_174 : L0Memory_45; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_275 = count >= 10'h1 & count <= _T_27 ? _GEN_175 : L0Memory_46; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_276 = count >= 10'h1 & count <= _T_27 ? _GEN_176 : L0Memory_47; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_277 = count >= 10'h1 & count <= _T_27 ? _GEN_177 : L0Memory_48; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_278 = count >= 10'h1 & count <= _T_27 ? _GEN_178 : L0Memory_49; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_279 = count >= 10'h1 & count <= _T_27 ? _GEN_179 : L0Memory_50; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_280 = count >= 10'h1 & count <= _T_27 ? _GEN_180 : L0Memory_51; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_281 = count >= 10'h1 & count <= _T_27 ? _GEN_181 : L0Memory_52; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_282 = count >= 10'h1 & count <= _T_27 ? _GEN_182 : L0Memory_53; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_283 = count >= 10'h1 & count <= _T_27 ? _GEN_183 : L0Memory_54; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_284 = count >= 10'h1 & count <= _T_27 ? _GEN_184 : L0Memory_55; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_285 = count >= 10'h1 & count <= _T_27 ? _GEN_185 : L0Memory_56; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_286 = count >= 10'h1 & count <= _T_27 ? _GEN_186 : L0Memory_57; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_287 = count >= 10'h1 & count <= _T_27 ? _GEN_187 : L0Memory_58; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_288 = count >= 10'h1 & count <= _T_27 ? _GEN_188 : L0Memory_59; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_289 = count >= 10'h1 & count <= _T_27 ? _GEN_189 : L0Memory_60; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_290 = count >= 10'h1 & count <= _T_27 ? _GEN_190 : L0Memory_61; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_291 = count >= 10'h1 & count <= _T_27 ? _GEN_191 : L0Memory_62; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_292 = count >= 10'h1 & count <= _T_27 ? _GEN_192 : L0Memory_63; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_293 = count >= 10'h1 & count <= _T_27 ? _GEN_193 : L0Memory_64; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_294 = count >= 10'h1 & count <= _T_27 ? _GEN_194 : L0Memory_65; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_295 = count >= 10'h1 & count <= _T_27 ? _GEN_195 : L0Memory_66; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_296 = count >= 10'h1 & count <= _T_27 ? _GEN_196 : L0Memory_67; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_297 = count >= 10'h1 & count <= _T_27 ? _GEN_197 : L0Memory_68; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_298 = count >= 10'h1 & count <= _T_27 ? _GEN_198 : L0Memory_69; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_299 = count >= 10'h1 & count <= _T_27 ? _GEN_199 : L0Memory_70; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_300 = count >= 10'h1 & count <= _T_27 ? _GEN_200 : L0Memory_71; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_301 = count >= 10'h1 & count <= _T_27 ? _GEN_201 : L0Memory_72; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_302 = count >= 10'h1 & count <= _T_27 ? _GEN_202 : L0Memory_73; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_303 = count >= 10'h1 & count <= _T_27 ? _GEN_203 : L0Memory_74; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_304 = count >= 10'h1 & count <= _T_27 ? _GEN_204 : L0Memory_75; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_305 = count >= 10'h1 & count <= _T_27 ? _GEN_205 : L0Memory_76; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_306 = count >= 10'h1 & count <= _T_27 ? _GEN_206 : L0Memory_77; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_307 = count >= 10'h1 & count <= _T_27 ? _GEN_207 : L0Memory_78; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_308 = count >= 10'h1 & count <= _T_27 ? _GEN_208 : L0Memory_79; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_309 = count >= 10'h1 & count <= _T_27 ? _GEN_209 : L0Memory_80; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_310 = count >= 10'h1 & count <= _T_27 ? _GEN_210 : L0Memory_81; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_311 = count >= 10'h1 & count <= _T_27 ? _GEN_211 : L0Memory_82; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_312 = count >= 10'h1 & count <= _T_27 ? _GEN_212 : L0Memory_83; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_313 = count >= 10'h1 & count <= _T_27 ? _GEN_213 : L0Memory_84; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_314 = count >= 10'h1 & count <= _T_27 ? _GEN_214 : L0Memory_85; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_315 = count >= 10'h1 & count <= _T_27 ? _GEN_215 : L0Memory_86; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_316 = count >= 10'h1 & count <= _T_27 ? _GEN_216 : L0Memory_87; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_317 = count >= 10'h1 & count <= _T_27 ? _GEN_217 : L0Memory_88; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_318 = count >= 10'h1 & count <= _T_27 ? _GEN_218 : L0Memory_89; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_319 = count >= 10'h1 & count <= _T_27 ? _GEN_219 : L0Memory_90; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_320 = count >= 10'h1 & count <= _T_27 ? _GEN_220 : L0Memory_91; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_321 = count >= 10'h1 & count <= _T_27 ? _GEN_221 : L0Memory_92; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_322 = count >= 10'h1 & count <= _T_27 ? _GEN_222 : L0Memory_93; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_323 = count >= 10'h1 & count <= _T_27 ? _GEN_223 : L0Memory_94; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_324 = count >= 10'h1 & count <= _T_27 ? _GEN_224 : L0Memory_95; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_325 = count >= 10'h1 & count <= _T_27 ? _GEN_225 : L0Memory_96; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_326 = count >= 10'h1 & count <= _T_27 ? _GEN_226 : L0Memory_97; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_327 = count >= 10'h1 & count <= _T_27 ? _GEN_227 : L0Memory_98; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_328 = count >= 10'h1 & count <= _T_27 ? _GEN_228 : L0Memory_99; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [5:0] _GEN_329 = count >= 10'h1 & count <= _T_27 ? _L0Index_T_2 : _GEN_128; // @[PEArray.scala 198:59 PEArray.scala 200:17]
  wire [9:0] _GEN_330 = _T_24 ? 10'h0 : _GEN_127; // @[PEArray.scala 202:32 PEArray.scala 203:15]
  wire [2:0] _GEN_331 = _T_24 ? 3'h0 : state; // @[PEArray.scala 202:32 PEArray.scala 204:15 PEArray.scala 100:22]
  wire [9:0] _GEN_865 = {{4'd0}, GRU_out_width}; // @[PEArray.scala 220:19]
  wire [9:0] _GEN_0 = count % _GEN_865; // @[PEArray.scala 220:19]
  wire [5:0] _T_36 = _GEN_0[5:0]; // @[PEArray.scala 220:19]
  wire [5:0] _T_38 = GRU_out_width - 6'h1; // @[PEArray.scala 220:55]
  wire [5:0] _GEN_334 = _T_36 == _T_38 ? _L0Index_T_2 : 6'h0; // @[PEArray.scala 220:62 PEArray.scala 221:17 PEArray.scala 214:15]
  wire [5:0] _GEN_346 = _T_41 ? _GEN_334 : L0Index; // @[Conditional.scala 39:67 PEArray.scala 39:24]
  wire [9:0] _GEN_347 = _T_41 ? _GEN_330 : count; // @[Conditional.scala 39:67 PEArray.scala 101:22]
  wire [2:0] _GEN_348 = _T_41 ? _GEN_331 : state; // @[Conditional.scala 39:67 PEArray.scala 100:22]
  wire [5:0] _GEN_353 = _T_31 ? _GEN_334 : _GEN_346; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_354 = _T_31 ? _GEN_330 : _GEN_347; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_355 = _T_31 ? _GEN_331 : _GEN_348; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_356 = _T_22 ? _GEN_330 : _GEN_354; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_357 = _T_22 ? _GEN_329 : _GEN_353; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_458 = _T_22 ? _GEN_331 : _GEN_355; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_690 = _T_3 ? _GEN_118 : {{2'd0}, GRU_out_width}; // @[Conditional.scala 40:58 PEArray.scala 104:26]
  FP16MulAdder FP16MAC ( // @[PEArray.scala 72:23]
    .io_a(FP16MAC_io_a),
    .io_b(FP16MAC_io_b),
    .io_c(FP16MAC_io_c),
    .io_out(FP16MAC_io_out)
  );
  assign io_ToRightPE = mux3out_reg; // @[PEArray.scala 95:16]
  assign io_ToBelowPE = mux2out_reg; // @[PEArray.scala 94:16]
  assign FP16MAC_io_a = sel1 ? io_FromL1 : io_FromLeftPE; // @[PEArray.scala 50:14 PEArray.scala 50:23 PEArray.scala 51:24]
  assign FP16MAC_io_b = sel5 ? mux4out : _GEN_105; // @[PEArray.scala 77:13 PEArray.scala 78:18 PEArray.scala 81:18]
  assign FP16MAC_io_c = sel5 ? _GEN_105 : mux4out; // @[PEArray.scala 77:13 PEArray.scala 79:18 PEArray.scala 82:18]
  always @(posedge clock) begin
    if (reset) begin // @[PEArray.scala 39:24]
      L0Index <= 6'h0; // @[PEArray.scala 39:24]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h1; // @[PEArray.scala 159:15]
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h4; // @[PEArray.scala 181:15]
      end else begin
        L0Index <= _GEN_357;
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_0 <= _GEN_229;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_1 <= _GEN_230;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_2 <= _GEN_231;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_3 <= _GEN_232;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_4 <= _GEN_233;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_5 <= _GEN_234;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_6 <= _GEN_235;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_7 <= _GEN_236;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_8 <= _GEN_237;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_9 <= _GEN_238;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_10 <= _GEN_239;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_11 <= _GEN_240;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_12 <= _GEN_241;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_13 <= _GEN_242;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_14 <= _GEN_243;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_15 <= _GEN_244;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_16 <= _GEN_245;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_17 <= _GEN_246;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_18 <= _GEN_247;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_19 <= _GEN_248;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_20 <= _GEN_249;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_21 <= _GEN_250;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_22 <= _GEN_251;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_23 <= _GEN_252;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_24 <= _GEN_253;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_25 <= _GEN_254;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_26 <= _GEN_255;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_27 <= _GEN_256;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_28 <= _GEN_257;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_29 <= _GEN_258;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_30 <= _GEN_259;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_31 <= _GEN_260;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_32 <= _GEN_261;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_33 <= _GEN_262;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_34 <= _GEN_263;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_35 <= _GEN_264;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_36 <= _GEN_265;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_37 <= _GEN_266;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_38 <= _GEN_267;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_39 <= _GEN_268;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_40 <= _GEN_269;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_41 <= _GEN_270;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_42 <= _GEN_271;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_43 <= _GEN_272;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_44 <= _GEN_273;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_45 <= _GEN_274;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_46 <= _GEN_275;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_47 <= _GEN_276;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_48 <= _GEN_277;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_49 <= _GEN_278;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_50 <= _GEN_279;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_51 <= _GEN_280;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_52 <= _GEN_281;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_53 <= _GEN_282;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_54 <= _GEN_283;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_55 <= _GEN_284;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_56 <= _GEN_285;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_57 <= _GEN_286;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_58 <= _GEN_287;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_59 <= _GEN_288;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_60 <= _GEN_289;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_61 <= _GEN_290;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_62 <= _GEN_291;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_63 <= _GEN_292;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_64 <= _GEN_293;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_65 <= _GEN_294;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_66 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_67 <= _GEN_296;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_68 <= _GEN_297;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_69 <= _GEN_298;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_70 <= _GEN_299;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_71 <= _GEN_300;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_72 <= _GEN_301;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_73 <= _GEN_302;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_74 <= _GEN_303;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_75 <= _GEN_304;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_76 <= _GEN_305;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_77 <= _GEN_306;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_78 <= _GEN_307;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_79 <= _GEN_308;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_80 <= _GEN_309;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_81 <= _GEN_310;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_82 <= _GEN_311;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_83 <= _GEN_312;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_84 <= _GEN_313;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_85 <= _GEN_314;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_86 <= _GEN_315;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_87 <= _GEN_316;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_88 <= _GEN_317;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_89 <= _GEN_318;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_90 <= _GEN_319;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_91 <= _GEN_320;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_92 <= _GEN_321;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_93 <= _GEN_322;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_94 <= _GEN_323;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_95 <= _GEN_324;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_96 <= _GEN_325;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_97 <= _GEN_326;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_98 <= _GEN_327;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_99 <= _GEN_328;
          end
        end
      end
    end
    if (reset) begin // @[PEArray.scala 100:22]
      state <= 3'h0; // @[PEArray.scala 100:22]
    end else if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[10]) begin // @[PEArray.scala 116:57]
        state <= 3'h1;
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      if (count == 10'h33) begin // @[PEArray.scala 164:27]
        state <= 3'h0; // @[PEArray.scala 166:15]
      end
    end else if (_T_16) begin // @[Conditional.scala 39:67]
      state <= _GEN_126;
    end else begin
      state <= _GEN_458;
    end
    if (reset) begin // @[PEArray.scala 90:28]
      mux2out_reg <= 16'h0; // @[PEArray.scala 90:28]
    end else begin
      mux2out_reg <= MAC_out; // @[PEArray.scala 90:28]
    end
    if (reset) begin // @[PEArray.scala 91:28]
      mux3out_reg <= 16'h0; // @[PEArray.scala 91:28]
    end else if (sel3) begin // @[PEArray.scala 56:14]
      mux3out_reg <= MAC_out; // @[PEArray.scala 56:23]
    end else if (sel1) begin // @[PEArray.scala 50:14]
      mux3out_reg <= io_FromL1; // @[PEArray.scala 50:23]
    end else begin
      mux3out_reg <= io_FromLeftPE; // @[PEArray.scala 51:24]
    end
    if (reset) begin // @[PEArray.scala 101:22]
      count <= 10'h0; // @[PEArray.scala 101:22]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        if (count == 10'h33) begin // @[PEArray.scala 164:27]
          count <= 10'h0; // @[PEArray.scala 165:15]
        end else begin
          count <= _GEN_120;
        end
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        count <= _GEN_125;
      end else begin
        count <= _GEN_356;
      end
    end
    GRU_out_width <= _GEN_690[5:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  L0Index = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  L0Memory_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  L0Memory_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  L0Memory_2 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  L0Memory_3 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  L0Memory_4 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  L0Memory_5 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  L0Memory_6 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  L0Memory_7 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  L0Memory_8 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  L0Memory_9 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  L0Memory_10 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  L0Memory_11 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  L0Memory_12 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  L0Memory_13 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  L0Memory_14 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  L0Memory_15 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  L0Memory_16 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  L0Memory_17 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  L0Memory_18 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  L0Memory_19 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  L0Memory_20 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  L0Memory_21 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  L0Memory_22 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  L0Memory_23 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  L0Memory_24 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  L0Memory_25 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  L0Memory_26 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  L0Memory_27 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  L0Memory_28 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  L0Memory_29 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  L0Memory_30 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  L0Memory_31 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  L0Memory_32 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  L0Memory_33 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  L0Memory_34 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  L0Memory_35 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  L0Memory_36 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  L0Memory_37 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  L0Memory_38 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  L0Memory_39 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  L0Memory_40 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  L0Memory_41 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  L0Memory_42 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  L0Memory_43 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  L0Memory_44 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  L0Memory_45 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  L0Memory_46 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  L0Memory_47 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  L0Memory_48 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  L0Memory_49 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  L0Memory_50 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  L0Memory_51 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  L0Memory_52 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  L0Memory_53 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  L0Memory_54 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  L0Memory_55 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  L0Memory_56 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  L0Memory_57 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  L0Memory_58 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  L0Memory_59 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  L0Memory_60 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  L0Memory_61 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  L0Memory_62 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  L0Memory_63 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  L0Memory_64 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  L0Memory_65 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  L0Memory_66 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  L0Memory_67 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  L0Memory_68 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  L0Memory_69 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  L0Memory_70 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  L0Memory_71 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  L0Memory_72 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  L0Memory_73 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  L0Memory_74 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  L0Memory_75 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  L0Memory_76 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  L0Memory_77 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  L0Memory_78 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  L0Memory_79 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  L0Memory_80 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  L0Memory_81 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  L0Memory_82 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  L0Memory_83 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  L0Memory_84 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  L0Memory_85 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  L0Memory_86 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  L0Memory_87 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  L0Memory_88 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  L0Memory_89 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  L0Memory_90 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  L0Memory_91 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  L0Memory_92 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  L0Memory_93 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  L0Memory_94 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  L0Memory_95 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  L0Memory_96 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  L0Memory_97 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  L0Memory_98 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  L0Memory_99 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  state = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  mux2out_reg = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  mux3out_reg = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  count = _RAND_104[9:0];
  _RAND_105 = {1{`RANDOM}};
  GRU_out_width = _RAND_105[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PE_5(
  input         clock,
  input         reset,
  input  [15:0] io_FromAbovePE,
  input  [15:0] io_FromLeftPE,
  input  [15:0] io_FromL1,
  input  [2:0]  io_control_signal_control,
  input  [9:0]  io_control_signal_count,
  input  [5:0]  io_control_signal_L0index,
  input  [11:0] io_control_signal_mask,
  input  [7:0]  io_control_signal_gru_out_width,
  output [15:0] io_ToRightPE,
  output [15:0] io_ToBelowPE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] FP16MAC_io_a; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_b; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_c; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_out; // @[PEArray.scala 72:23]
  reg [5:0] L0Index; // @[PEArray.scala 39:24]
  reg [15:0] L0Memory_0; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_1; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_2; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_3; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_4; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_5; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_6; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_7; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_8; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_9; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_10; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_11; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_12; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_13; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_14; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_15; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_16; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_17; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_18; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_19; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_20; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_21; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_22; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_23; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_24; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_25; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_26; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_27; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_28; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_29; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_30; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_31; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_32; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_33; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_34; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_35; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_36; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_37; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_38; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_39; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_40; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_41; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_42; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_43; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_44; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_45; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_46; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_47; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_48; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_49; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_50; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_51; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_52; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_53; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_54; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_55; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_56; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_57; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_58; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_59; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_60; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_61; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_62; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_63; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_64; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_65; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_66; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_67; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_68; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_69; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_70; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_71; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_72; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_73; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_74; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_75; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_76; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_77; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_78; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_79; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_80; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_81; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_82; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_83; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_84; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_85; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_86; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_87; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_88; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_89; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_90; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_91; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_92; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_93; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_94; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_95; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_96; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_97; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_98; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_99; // @[PEArray.scala 40:21]
  reg [2:0] state; // @[PEArray.scala 100:22]
  wire  _T_3 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_12 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_16 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_22 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_31 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_41 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_342 = _T_41 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 231:12 PEArray.scala 32:8]
  wire  _GEN_349 = _T_31 ? 1'h0 : _GEN_342; // @[Conditional.scala 39:67 PEArray.scala 208:12]
  wire  _GEN_459 = _T_22 | _GEN_349; // @[Conditional.scala 39:67 PEArray.scala 32:8]
  wire  _GEN_463 = _T_16 ? 1'h0 : _GEN_459; // @[Conditional.scala 39:67]
  wire  _GEN_572 = _T_12 | _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 149:12]
  wire  sel1 = _T_3 | _GEN_572; // @[Conditional.scala 40:58 PEArray.scala 108:12]
  wire [15:0] MAC_out = FP16MAC_io_out; // @[PEArray.scala 47:21 PEArray.scala 85:11]
  wire  _GEN_465 = _T_16 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 177:12]
  wire  _GEN_580 = _T_12 | _GEN_465; // @[Conditional.scala 39:67 PEArray.scala 34:8]
  wire  sel3 = _T_3 | _GEN_580; // @[Conditional.scala 40:58 PEArray.scala 110:12]
  wire [1:0] _GEN_344 = _T_41 ? 2'h2 : 2'h0; // @[Conditional.scala 39:67 PEArray.scala 233:12 PEArray.scala 35:8]
  wire [1:0] _GEN_351 = _T_31 ? 2'h2 : _GEN_344; // @[Conditional.scala 39:67 PEArray.scala 210:12]
  wire [1:0] _GEN_461 = _T_22 ? 2'h0 : _GEN_351; // @[Conditional.scala 39:67 PEArray.scala 35:8]
  wire [1:0] _GEN_466 = _T_16 ? 2'h0 : _GEN_461; // @[Conditional.scala 39:67 PEArray.scala 178:12]
  wire [1:0] _GEN_574 = _T_12 ? 2'h1 : _GEN_466; // @[Conditional.scala 39:67]
  wire [1:0] sel4 = _T_3 ? 2'h0 : _GEN_574; // @[Conditional.scala 40:58 PEArray.scala 111:12]
  wire [15:0] _GEN_3 = sel4 == 2'h2 ? io_FromL1 : 16'h0; // @[PEArray.scala 65:28 PEArray.scala 66:15 PEArray.scala 69:15]
  wire [15:0] _GEN_4 = sel4 == 2'h1 ? io_FromAbovePE : _GEN_3; // @[PEArray.scala 62:28 PEArray.scala 63:15]
  wire [15:0] mux4out = sel4 == 2'h0 ? 16'h0 : _GEN_4; // @[PEArray.scala 59:22 PEArray.scala 60:13]
  wire [15:0] _GEN_7 = 6'h1 == L0Index ? L0Memory_1 : L0Memory_0; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_8 = 6'h2 == L0Index ? L0Memory_2 : _GEN_7; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_9 = 6'h3 == L0Index ? L0Memory_3 : _GEN_8; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_10 = 6'h4 == L0Index ? L0Memory_4 : _GEN_9; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_11 = 6'h5 == L0Index ? L0Memory_5 : _GEN_10; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_12 = 6'h6 == L0Index ? L0Memory_6 : _GEN_11; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_13 = 6'h7 == L0Index ? L0Memory_7 : _GEN_12; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_14 = 6'h8 == L0Index ? L0Memory_8 : _GEN_13; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_15 = 6'h9 == L0Index ? L0Memory_9 : _GEN_14; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_16 = 6'ha == L0Index ? L0Memory_10 : _GEN_15; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_17 = 6'hb == L0Index ? L0Memory_11 : _GEN_16; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_18 = 6'hc == L0Index ? L0Memory_12 : _GEN_17; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_19 = 6'hd == L0Index ? L0Memory_13 : _GEN_18; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_20 = 6'he == L0Index ? L0Memory_14 : _GEN_19; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_21 = 6'hf == L0Index ? L0Memory_15 : _GEN_20; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_22 = 6'h10 == L0Index ? L0Memory_16 : _GEN_21; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_23 = 6'h11 == L0Index ? L0Memory_17 : _GEN_22; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_24 = 6'h12 == L0Index ? L0Memory_18 : _GEN_23; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_25 = 6'h13 == L0Index ? L0Memory_19 : _GEN_24; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_26 = 6'h14 == L0Index ? L0Memory_20 : _GEN_25; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_27 = 6'h15 == L0Index ? L0Memory_21 : _GEN_26; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_28 = 6'h16 == L0Index ? L0Memory_22 : _GEN_27; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_29 = 6'h17 == L0Index ? L0Memory_23 : _GEN_28; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_30 = 6'h18 == L0Index ? L0Memory_24 : _GEN_29; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_31 = 6'h19 == L0Index ? L0Memory_25 : _GEN_30; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_32 = 6'h1a == L0Index ? L0Memory_26 : _GEN_31; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_33 = 6'h1b == L0Index ? L0Memory_27 : _GEN_32; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_34 = 6'h1c == L0Index ? L0Memory_28 : _GEN_33; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_35 = 6'h1d == L0Index ? L0Memory_29 : _GEN_34; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_36 = 6'h1e == L0Index ? L0Memory_30 : _GEN_35; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_37 = 6'h1f == L0Index ? L0Memory_31 : _GEN_36; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_38 = 6'h20 == L0Index ? L0Memory_32 : _GEN_37; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_39 = 6'h21 == L0Index ? L0Memory_33 : _GEN_38; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_40 = 6'h22 == L0Index ? L0Memory_34 : _GEN_39; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_41 = 6'h23 == L0Index ? L0Memory_35 : _GEN_40; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_42 = 6'h24 == L0Index ? L0Memory_36 : _GEN_41; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_43 = 6'h25 == L0Index ? L0Memory_37 : _GEN_42; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_44 = 6'h26 == L0Index ? L0Memory_38 : _GEN_43; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_45 = 6'h27 == L0Index ? L0Memory_39 : _GEN_44; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_46 = 6'h28 == L0Index ? L0Memory_40 : _GEN_45; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_47 = 6'h29 == L0Index ? L0Memory_41 : _GEN_46; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_48 = 6'h2a == L0Index ? L0Memory_42 : _GEN_47; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_49 = 6'h2b == L0Index ? L0Memory_43 : _GEN_48; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_50 = 6'h2c == L0Index ? L0Memory_44 : _GEN_49; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_51 = 6'h2d == L0Index ? L0Memory_45 : _GEN_50; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_52 = 6'h2e == L0Index ? L0Memory_46 : _GEN_51; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_53 = 6'h2f == L0Index ? L0Memory_47 : _GEN_52; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_54 = 6'h30 == L0Index ? L0Memory_48 : _GEN_53; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_55 = 6'h31 == L0Index ? L0Memory_49 : _GEN_54; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_56 = 6'h32 == L0Index ? L0Memory_50 : _GEN_55; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_57 = 6'h33 == L0Index ? L0Memory_51 : _GEN_56; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_58 = 6'h34 == L0Index ? L0Memory_52 : _GEN_57; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_59 = 6'h35 == L0Index ? L0Memory_53 : _GEN_58; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_60 = 6'h36 == L0Index ? L0Memory_54 : _GEN_59; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_61 = 6'h37 == L0Index ? L0Memory_55 : _GEN_60; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_62 = 6'h38 == L0Index ? L0Memory_56 : _GEN_61; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_63 = 6'h39 == L0Index ? L0Memory_57 : _GEN_62; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_64 = 6'h3a == L0Index ? L0Memory_58 : _GEN_63; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_65 = 6'h3b == L0Index ? L0Memory_59 : _GEN_64; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_66 = 6'h3c == L0Index ? L0Memory_60 : _GEN_65; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_67 = 6'h3d == L0Index ? L0Memory_61 : _GEN_66; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_68 = 6'h3e == L0Index ? L0Memory_62 : _GEN_67; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_69 = 6'h3f == L0Index ? L0Memory_63 : _GEN_68; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [6:0] _GEN_793 = {{1'd0}, L0Index}; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_70 = 7'h40 == _GEN_793 ? L0Memory_64 : _GEN_69; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_71 = 7'h41 == _GEN_793 ? L0Memory_65 : _GEN_70; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_72 = 7'h42 == _GEN_793 ? L0Memory_66 : _GEN_71; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_73 = 7'h43 == _GEN_793 ? L0Memory_67 : _GEN_72; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_74 = 7'h44 == _GEN_793 ? L0Memory_68 : _GEN_73; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_75 = 7'h45 == _GEN_793 ? L0Memory_69 : _GEN_74; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_76 = 7'h46 == _GEN_793 ? L0Memory_70 : _GEN_75; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_77 = 7'h47 == _GEN_793 ? L0Memory_71 : _GEN_76; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_78 = 7'h48 == _GEN_793 ? L0Memory_72 : _GEN_77; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_79 = 7'h49 == _GEN_793 ? L0Memory_73 : _GEN_78; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_80 = 7'h4a == _GEN_793 ? L0Memory_74 : _GEN_79; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_81 = 7'h4b == _GEN_793 ? L0Memory_75 : _GEN_80; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_82 = 7'h4c == _GEN_793 ? L0Memory_76 : _GEN_81; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_83 = 7'h4d == _GEN_793 ? L0Memory_77 : _GEN_82; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_84 = 7'h4e == _GEN_793 ? L0Memory_78 : _GEN_83; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_85 = 7'h4f == _GEN_793 ? L0Memory_79 : _GEN_84; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_86 = 7'h50 == _GEN_793 ? L0Memory_80 : _GEN_85; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_87 = 7'h51 == _GEN_793 ? L0Memory_81 : _GEN_86; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_88 = 7'h52 == _GEN_793 ? L0Memory_82 : _GEN_87; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_89 = 7'h53 == _GEN_793 ? L0Memory_83 : _GEN_88; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_90 = 7'h54 == _GEN_793 ? L0Memory_84 : _GEN_89; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_91 = 7'h55 == _GEN_793 ? L0Memory_85 : _GEN_90; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_92 = 7'h56 == _GEN_793 ? L0Memory_86 : _GEN_91; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_93 = 7'h57 == _GEN_793 ? L0Memory_87 : _GEN_92; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_94 = 7'h58 == _GEN_793 ? L0Memory_88 : _GEN_93; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_95 = 7'h59 == _GEN_793 ? L0Memory_89 : _GEN_94; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_96 = 7'h5a == _GEN_793 ? L0Memory_90 : _GEN_95; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_97 = 7'h5b == _GEN_793 ? L0Memory_91 : _GEN_96; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_98 = 7'h5c == _GEN_793 ? L0Memory_92 : _GEN_97; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_99 = 7'h5d == _GEN_793 ? L0Memory_93 : _GEN_98; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_100 = 7'h5e == _GEN_793 ? L0Memory_94 : _GEN_99; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_101 = 7'h5f == _GEN_793 ? L0Memory_95 : _GEN_100; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_102 = 7'h60 == _GEN_793 ? L0Memory_96 : _GEN_101; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_103 = 7'h61 == _GEN_793 ? L0Memory_97 : _GEN_102; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_104 = 7'h62 == _GEN_793 ? L0Memory_98 : _GEN_103; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_105 = 7'h63 == _GEN_793 ? L0Memory_99 : _GEN_104; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire  _GEN_575 = _T_12 ? 1'h0 : _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 157:12]
  wire  sel5 = _T_3 ? 1'h0 : _GEN_575; // @[Conditional.scala 40:58 PEArray.scala 112:12]
  reg [15:0] mux2out_reg; // @[PEArray.scala 90:28]
  reg [15:0] mux3out_reg; // @[PEArray.scala 91:28]
  reg [9:0] count; // @[PEArray.scala 101:22]
  reg [9:0] count_max; // @[PEArray.scala 102:22]
  reg [5:0] L0index_begin; // @[PEArray.scala 103:26]
  reg [5:0] GRU_out_width; // @[PEArray.scala 104:26]
  wire  _T_6 = 3'h0 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_7 = 3'h1 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_8 = 3'h2 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_9 = 3'h3 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_10 = 3'h4 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_11 = 3'h5 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_109 = _T_11 ? 3'h5 : state; // @[Conditional.scala 39:67 PEArray.scala 140:19 PEArray.scala 100:22]
  wire [2:0] _GEN_110 = _T_10 ? 3'h4 : _GEN_109; // @[Conditional.scala 39:67 PEArray.scala 136:19]
  wire [2:0] _GEN_111 = _T_9 ? 3'h3 : _GEN_110; // @[Conditional.scala 39:67 PEArray.scala 132:19]
  wire [2:0] _GEN_112 = _T_8 ? 3'h2 : _GEN_111; // @[Conditional.scala 39:67 PEArray.scala 128:19]
  wire [2:0] _GEN_113 = _T_7 ? 3'h1 : _GEN_112; // @[Conditional.scala 39:67 PEArray.scala 124:19]
  wire [7:0] _GEN_118 = io_control_signal_mask[10] ? io_control_signal_gru_out_width : {{2'd0}, GRU_out_width}; // @[PEArray.scala 116:57 PEArray.scala 145:23 PEArray.scala 104:26]
  wire [9:0] _count_T_1 = count + 10'h1; // @[PEArray.scala 162:24]
  wire [9:0] _GEN_120 = count != 10'h33 ? _count_T_1 : count; // @[PEArray.scala 161:27 PEArray.scala 162:15 PEArray.scala 101:22]
  wire [9:0] _GEN_124 = count != 10'h188 ? _count_T_1 : count; // @[PEArray.scala 183:28 PEArray.scala 184:15 PEArray.scala 101:22]
  wire [9:0] _GEN_125 = count == 10'h188 ? 10'h0 : _GEN_124; // @[PEArray.scala 186:28 PEArray.scala 187:15]
  wire [2:0] _GEN_126 = count == 10'h188 ? 3'h0 : state; // @[PEArray.scala 186:28 PEArray.scala 188:15 PEArray.scala 100:22]
  wire [9:0] _GEN_127 = count != count_max ? _count_T_1 : count; // @[PEArray.scala 192:32 PEArray.scala 193:15 PEArray.scala 101:22]
  wire [5:0] _GEN_128 = count == 10'h0 ? L0index_begin : L0Index; // @[PEArray.scala 195:26 PEArray.scala 196:17 PEArray.scala 39:24]
  wire [9:0] _T_27 = count_max - 10'h1; // @[PEArray.scala 198:51]
  wire [15:0] _GEN_129 = 6'h0 == L0Index ? io_FromL1 : L0Memory_0; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_130 = 6'h1 == L0Index ? io_FromL1 : L0Memory_1; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_131 = 6'h2 == L0Index ? io_FromL1 : L0Memory_2; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_132 = 6'h3 == L0Index ? io_FromL1 : L0Memory_3; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_133 = 6'h4 == L0Index ? io_FromL1 : L0Memory_4; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_134 = 6'h5 == L0Index ? io_FromL1 : L0Memory_5; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_135 = 6'h6 == L0Index ? io_FromL1 : L0Memory_6; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_136 = 6'h7 == L0Index ? io_FromL1 : L0Memory_7; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_137 = 6'h8 == L0Index ? io_FromL1 : L0Memory_8; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_138 = 6'h9 == L0Index ? io_FromL1 : L0Memory_9; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_139 = 6'ha == L0Index ? io_FromL1 : L0Memory_10; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_140 = 6'hb == L0Index ? io_FromL1 : L0Memory_11; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_141 = 6'hc == L0Index ? io_FromL1 : L0Memory_12; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_142 = 6'hd == L0Index ? io_FromL1 : L0Memory_13; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_143 = 6'he == L0Index ? io_FromL1 : L0Memory_14; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_144 = 6'hf == L0Index ? io_FromL1 : L0Memory_15; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_145 = 6'h10 == L0Index ? io_FromL1 : L0Memory_16; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_146 = 6'h11 == L0Index ? io_FromL1 : L0Memory_17; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_147 = 6'h12 == L0Index ? io_FromL1 : L0Memory_18; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_148 = 6'h13 == L0Index ? io_FromL1 : L0Memory_19; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_149 = 6'h14 == L0Index ? io_FromL1 : L0Memory_20; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_150 = 6'h15 == L0Index ? io_FromL1 : L0Memory_21; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_151 = 6'h16 == L0Index ? io_FromL1 : L0Memory_22; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_152 = 6'h17 == L0Index ? io_FromL1 : L0Memory_23; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_153 = 6'h18 == L0Index ? io_FromL1 : L0Memory_24; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_154 = 6'h19 == L0Index ? io_FromL1 : L0Memory_25; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_155 = 6'h1a == L0Index ? io_FromL1 : L0Memory_26; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_156 = 6'h1b == L0Index ? io_FromL1 : L0Memory_27; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_157 = 6'h1c == L0Index ? io_FromL1 : L0Memory_28; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_158 = 6'h1d == L0Index ? io_FromL1 : L0Memory_29; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_159 = 6'h1e == L0Index ? io_FromL1 : L0Memory_30; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_160 = 6'h1f == L0Index ? io_FromL1 : L0Memory_31; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_161 = 6'h20 == L0Index ? io_FromL1 : L0Memory_32; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_162 = 6'h21 == L0Index ? io_FromL1 : L0Memory_33; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_163 = 6'h22 == L0Index ? io_FromL1 : L0Memory_34; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_164 = 6'h23 == L0Index ? io_FromL1 : L0Memory_35; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_165 = 6'h24 == L0Index ? io_FromL1 : L0Memory_36; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_166 = 6'h25 == L0Index ? io_FromL1 : L0Memory_37; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_167 = 6'h26 == L0Index ? io_FromL1 : L0Memory_38; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_168 = 6'h27 == L0Index ? io_FromL1 : L0Memory_39; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_169 = 6'h28 == L0Index ? io_FromL1 : L0Memory_40; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_170 = 6'h29 == L0Index ? io_FromL1 : L0Memory_41; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_171 = 6'h2a == L0Index ? io_FromL1 : L0Memory_42; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_172 = 6'h2b == L0Index ? io_FromL1 : L0Memory_43; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_173 = 6'h2c == L0Index ? io_FromL1 : L0Memory_44; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_174 = 6'h2d == L0Index ? io_FromL1 : L0Memory_45; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_175 = 6'h2e == L0Index ? io_FromL1 : L0Memory_46; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_176 = 6'h2f == L0Index ? io_FromL1 : L0Memory_47; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_177 = 6'h30 == L0Index ? io_FromL1 : L0Memory_48; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_178 = 6'h31 == L0Index ? io_FromL1 : L0Memory_49; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_179 = 6'h32 == L0Index ? io_FromL1 : L0Memory_50; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_180 = 6'h33 == L0Index ? io_FromL1 : L0Memory_51; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_181 = 6'h34 == L0Index ? io_FromL1 : L0Memory_52; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_182 = 6'h35 == L0Index ? io_FromL1 : L0Memory_53; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_183 = 6'h36 == L0Index ? io_FromL1 : L0Memory_54; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_184 = 6'h37 == L0Index ? io_FromL1 : L0Memory_55; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_185 = 6'h38 == L0Index ? io_FromL1 : L0Memory_56; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_186 = 6'h39 == L0Index ? io_FromL1 : L0Memory_57; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_187 = 6'h3a == L0Index ? io_FromL1 : L0Memory_58; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_188 = 6'h3b == L0Index ? io_FromL1 : L0Memory_59; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_189 = 6'h3c == L0Index ? io_FromL1 : L0Memory_60; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_190 = 6'h3d == L0Index ? io_FromL1 : L0Memory_61; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_191 = 6'h3e == L0Index ? io_FromL1 : L0Memory_62; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_192 = 6'h3f == L0Index ? io_FromL1 : L0Memory_63; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_193 = 7'h40 == _GEN_793 ? io_FromL1 : L0Memory_64; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_194 = 7'h41 == _GEN_793 ? io_FromL1 : L0Memory_65; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_195 = 7'h42 == _GEN_793 ? io_FromL1 : L0Memory_66; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_196 = 7'h43 == _GEN_793 ? io_FromL1 : L0Memory_67; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_197 = 7'h44 == _GEN_793 ? io_FromL1 : L0Memory_68; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_198 = 7'h45 == _GEN_793 ? io_FromL1 : L0Memory_69; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_199 = 7'h46 == _GEN_793 ? io_FromL1 : L0Memory_70; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_200 = 7'h47 == _GEN_793 ? io_FromL1 : L0Memory_71; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_201 = 7'h48 == _GEN_793 ? io_FromL1 : L0Memory_72; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_202 = 7'h49 == _GEN_793 ? io_FromL1 : L0Memory_73; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_203 = 7'h4a == _GEN_793 ? io_FromL1 : L0Memory_74; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_204 = 7'h4b == _GEN_793 ? io_FromL1 : L0Memory_75; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_205 = 7'h4c == _GEN_793 ? io_FromL1 : L0Memory_76; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_206 = 7'h4d == _GEN_793 ? io_FromL1 : L0Memory_77; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_207 = 7'h4e == _GEN_793 ? io_FromL1 : L0Memory_78; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_208 = 7'h4f == _GEN_793 ? io_FromL1 : L0Memory_79; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_209 = 7'h50 == _GEN_793 ? io_FromL1 : L0Memory_80; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_210 = 7'h51 == _GEN_793 ? io_FromL1 : L0Memory_81; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_211 = 7'h52 == _GEN_793 ? io_FromL1 : L0Memory_82; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_212 = 7'h53 == _GEN_793 ? io_FromL1 : L0Memory_83; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_213 = 7'h54 == _GEN_793 ? io_FromL1 : L0Memory_84; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_214 = 7'h55 == _GEN_793 ? io_FromL1 : L0Memory_85; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_215 = 7'h56 == _GEN_793 ? io_FromL1 : L0Memory_86; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_216 = 7'h57 == _GEN_793 ? io_FromL1 : L0Memory_87; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_217 = 7'h58 == _GEN_793 ? io_FromL1 : L0Memory_88; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_218 = 7'h59 == _GEN_793 ? io_FromL1 : L0Memory_89; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_219 = 7'h5a == _GEN_793 ? io_FromL1 : L0Memory_90; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_220 = 7'h5b == _GEN_793 ? io_FromL1 : L0Memory_91; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_221 = 7'h5c == _GEN_793 ? io_FromL1 : L0Memory_92; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_222 = 7'h5d == _GEN_793 ? io_FromL1 : L0Memory_93; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_223 = 7'h5e == _GEN_793 ? io_FromL1 : L0Memory_94; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_224 = 7'h5f == _GEN_793 ? io_FromL1 : L0Memory_95; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_225 = 7'h60 == _GEN_793 ? io_FromL1 : L0Memory_96; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_226 = 7'h61 == _GEN_793 ? io_FromL1 : L0Memory_97; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_227 = 7'h62 == _GEN_793 ? io_FromL1 : L0Memory_98; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_228 = 7'h63 == _GEN_793 ? io_FromL1 : L0Memory_99; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [5:0] _L0Index_T_2 = L0Index + 6'h1; // @[PEArray.scala 200:28]
  wire [15:0] _GEN_229 = count >= 10'h1 & count <= _T_27 ? _GEN_129 : L0Memory_0; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_230 = count >= 10'h1 & count <= _T_27 ? _GEN_130 : L0Memory_1; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_231 = count >= 10'h1 & count <= _T_27 ? _GEN_131 : L0Memory_2; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_232 = count >= 10'h1 & count <= _T_27 ? _GEN_132 : L0Memory_3; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_233 = count >= 10'h1 & count <= _T_27 ? _GEN_133 : L0Memory_4; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_234 = count >= 10'h1 & count <= _T_27 ? _GEN_134 : L0Memory_5; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_235 = count >= 10'h1 & count <= _T_27 ? _GEN_135 : L0Memory_6; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_236 = count >= 10'h1 & count <= _T_27 ? _GEN_136 : L0Memory_7; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_237 = count >= 10'h1 & count <= _T_27 ? _GEN_137 : L0Memory_8; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_238 = count >= 10'h1 & count <= _T_27 ? _GEN_138 : L0Memory_9; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_239 = count >= 10'h1 & count <= _T_27 ? _GEN_139 : L0Memory_10; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_240 = count >= 10'h1 & count <= _T_27 ? _GEN_140 : L0Memory_11; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_241 = count >= 10'h1 & count <= _T_27 ? _GEN_141 : L0Memory_12; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_242 = count >= 10'h1 & count <= _T_27 ? _GEN_142 : L0Memory_13; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_243 = count >= 10'h1 & count <= _T_27 ? _GEN_143 : L0Memory_14; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_244 = count >= 10'h1 & count <= _T_27 ? _GEN_144 : L0Memory_15; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_245 = count >= 10'h1 & count <= _T_27 ? _GEN_145 : L0Memory_16; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_246 = count >= 10'h1 & count <= _T_27 ? _GEN_146 : L0Memory_17; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_247 = count >= 10'h1 & count <= _T_27 ? _GEN_147 : L0Memory_18; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_248 = count >= 10'h1 & count <= _T_27 ? _GEN_148 : L0Memory_19; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_249 = count >= 10'h1 & count <= _T_27 ? _GEN_149 : L0Memory_20; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_250 = count >= 10'h1 & count <= _T_27 ? _GEN_150 : L0Memory_21; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_251 = count >= 10'h1 & count <= _T_27 ? _GEN_151 : L0Memory_22; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_252 = count >= 10'h1 & count <= _T_27 ? _GEN_152 : L0Memory_23; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_253 = count >= 10'h1 & count <= _T_27 ? _GEN_153 : L0Memory_24; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_254 = count >= 10'h1 & count <= _T_27 ? _GEN_154 : L0Memory_25; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_255 = count >= 10'h1 & count <= _T_27 ? _GEN_155 : L0Memory_26; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_256 = count >= 10'h1 & count <= _T_27 ? _GEN_156 : L0Memory_27; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_257 = count >= 10'h1 & count <= _T_27 ? _GEN_157 : L0Memory_28; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_258 = count >= 10'h1 & count <= _T_27 ? _GEN_158 : L0Memory_29; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_259 = count >= 10'h1 & count <= _T_27 ? _GEN_159 : L0Memory_30; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_260 = count >= 10'h1 & count <= _T_27 ? _GEN_160 : L0Memory_31; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_261 = count >= 10'h1 & count <= _T_27 ? _GEN_161 : L0Memory_32; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_262 = count >= 10'h1 & count <= _T_27 ? _GEN_162 : L0Memory_33; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_263 = count >= 10'h1 & count <= _T_27 ? _GEN_163 : L0Memory_34; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_264 = count >= 10'h1 & count <= _T_27 ? _GEN_164 : L0Memory_35; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_265 = count >= 10'h1 & count <= _T_27 ? _GEN_165 : L0Memory_36; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_266 = count >= 10'h1 & count <= _T_27 ? _GEN_166 : L0Memory_37; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_267 = count >= 10'h1 & count <= _T_27 ? _GEN_167 : L0Memory_38; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_268 = count >= 10'h1 & count <= _T_27 ? _GEN_168 : L0Memory_39; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_269 = count >= 10'h1 & count <= _T_27 ? _GEN_169 : L0Memory_40; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_270 = count >= 10'h1 & count <= _T_27 ? _GEN_170 : L0Memory_41; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_271 = count >= 10'h1 & count <= _T_27 ? _GEN_171 : L0Memory_42; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_272 = count >= 10'h1 & count <= _T_27 ? _GEN_172 : L0Memory_43; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_273 = count >= 10'h1 & count <= _T_27 ? _GEN_173 : L0Memory_44; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_274 = count >= 10'h1 & count <= _T_27 ? _GEN_174 : L0Memory_45; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_275 = count >= 10'h1 & count <= _T_27 ? _GEN_175 : L0Memory_46; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_276 = count >= 10'h1 & count <= _T_27 ? _GEN_176 : L0Memory_47; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_277 = count >= 10'h1 & count <= _T_27 ? _GEN_177 : L0Memory_48; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_278 = count >= 10'h1 & count <= _T_27 ? _GEN_178 : L0Memory_49; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_279 = count >= 10'h1 & count <= _T_27 ? _GEN_179 : L0Memory_50; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_280 = count >= 10'h1 & count <= _T_27 ? _GEN_180 : L0Memory_51; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_281 = count >= 10'h1 & count <= _T_27 ? _GEN_181 : L0Memory_52; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_282 = count >= 10'h1 & count <= _T_27 ? _GEN_182 : L0Memory_53; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_283 = count >= 10'h1 & count <= _T_27 ? _GEN_183 : L0Memory_54; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_284 = count >= 10'h1 & count <= _T_27 ? _GEN_184 : L0Memory_55; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_285 = count >= 10'h1 & count <= _T_27 ? _GEN_185 : L0Memory_56; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_286 = count >= 10'h1 & count <= _T_27 ? _GEN_186 : L0Memory_57; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_287 = count >= 10'h1 & count <= _T_27 ? _GEN_187 : L0Memory_58; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_288 = count >= 10'h1 & count <= _T_27 ? _GEN_188 : L0Memory_59; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_289 = count >= 10'h1 & count <= _T_27 ? _GEN_189 : L0Memory_60; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_290 = count >= 10'h1 & count <= _T_27 ? _GEN_190 : L0Memory_61; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_291 = count >= 10'h1 & count <= _T_27 ? _GEN_191 : L0Memory_62; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_292 = count >= 10'h1 & count <= _T_27 ? _GEN_192 : L0Memory_63; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_293 = count >= 10'h1 & count <= _T_27 ? _GEN_193 : L0Memory_64; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_294 = count >= 10'h1 & count <= _T_27 ? _GEN_194 : L0Memory_65; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_295 = count >= 10'h1 & count <= _T_27 ? _GEN_195 : L0Memory_66; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_296 = count >= 10'h1 & count <= _T_27 ? _GEN_196 : L0Memory_67; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_297 = count >= 10'h1 & count <= _T_27 ? _GEN_197 : L0Memory_68; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_298 = count >= 10'h1 & count <= _T_27 ? _GEN_198 : L0Memory_69; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_299 = count >= 10'h1 & count <= _T_27 ? _GEN_199 : L0Memory_70; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_300 = count >= 10'h1 & count <= _T_27 ? _GEN_200 : L0Memory_71; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_301 = count >= 10'h1 & count <= _T_27 ? _GEN_201 : L0Memory_72; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_302 = count >= 10'h1 & count <= _T_27 ? _GEN_202 : L0Memory_73; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_303 = count >= 10'h1 & count <= _T_27 ? _GEN_203 : L0Memory_74; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_304 = count >= 10'h1 & count <= _T_27 ? _GEN_204 : L0Memory_75; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_305 = count >= 10'h1 & count <= _T_27 ? _GEN_205 : L0Memory_76; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_306 = count >= 10'h1 & count <= _T_27 ? _GEN_206 : L0Memory_77; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_307 = count >= 10'h1 & count <= _T_27 ? _GEN_207 : L0Memory_78; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_308 = count >= 10'h1 & count <= _T_27 ? _GEN_208 : L0Memory_79; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_309 = count >= 10'h1 & count <= _T_27 ? _GEN_209 : L0Memory_80; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_310 = count >= 10'h1 & count <= _T_27 ? _GEN_210 : L0Memory_81; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_311 = count >= 10'h1 & count <= _T_27 ? _GEN_211 : L0Memory_82; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_312 = count >= 10'h1 & count <= _T_27 ? _GEN_212 : L0Memory_83; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_313 = count >= 10'h1 & count <= _T_27 ? _GEN_213 : L0Memory_84; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_314 = count >= 10'h1 & count <= _T_27 ? _GEN_214 : L0Memory_85; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_315 = count >= 10'h1 & count <= _T_27 ? _GEN_215 : L0Memory_86; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_316 = count >= 10'h1 & count <= _T_27 ? _GEN_216 : L0Memory_87; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_317 = count >= 10'h1 & count <= _T_27 ? _GEN_217 : L0Memory_88; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_318 = count >= 10'h1 & count <= _T_27 ? _GEN_218 : L0Memory_89; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_319 = count >= 10'h1 & count <= _T_27 ? _GEN_219 : L0Memory_90; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_320 = count >= 10'h1 & count <= _T_27 ? _GEN_220 : L0Memory_91; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_321 = count >= 10'h1 & count <= _T_27 ? _GEN_221 : L0Memory_92; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_322 = count >= 10'h1 & count <= _T_27 ? _GEN_222 : L0Memory_93; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_323 = count >= 10'h1 & count <= _T_27 ? _GEN_223 : L0Memory_94; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_324 = count >= 10'h1 & count <= _T_27 ? _GEN_224 : L0Memory_95; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_325 = count >= 10'h1 & count <= _T_27 ? _GEN_225 : L0Memory_96; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_326 = count >= 10'h1 & count <= _T_27 ? _GEN_226 : L0Memory_97; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_327 = count >= 10'h1 & count <= _T_27 ? _GEN_227 : L0Memory_98; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_328 = count >= 10'h1 & count <= _T_27 ? _GEN_228 : L0Memory_99; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [5:0] _GEN_329 = count >= 10'h1 & count <= _T_27 ? _L0Index_T_2 : _GEN_128; // @[PEArray.scala 198:59 PEArray.scala 200:17]
  wire [9:0] _GEN_330 = count == count_max ? 10'h0 : _GEN_127; // @[PEArray.scala 202:32 PEArray.scala 203:15]
  wire [2:0] _GEN_331 = count == count_max ? 3'h0 : state; // @[PEArray.scala 202:32 PEArray.scala 204:15 PEArray.scala 100:22]
  wire [9:0] _GEN_865 = {{4'd0}, GRU_out_width}; // @[PEArray.scala 220:19]
  wire [9:0] _GEN_0 = count % _GEN_865; // @[PEArray.scala 220:19]
  wire [5:0] _T_36 = _GEN_0[5:0]; // @[PEArray.scala 220:19]
  wire [5:0] _T_38 = GRU_out_width - 6'h1; // @[PEArray.scala 220:55]
  wire [5:0] _GEN_334 = _T_36 == _T_38 ? _L0Index_T_2 : L0index_begin; // @[PEArray.scala 220:62 PEArray.scala 221:17 PEArray.scala 214:15]
  wire [5:0] _GEN_346 = _T_41 ? _GEN_334 : L0Index; // @[Conditional.scala 39:67 PEArray.scala 39:24]
  wire [9:0] _GEN_347 = _T_41 ? _GEN_330 : count; // @[Conditional.scala 39:67 PEArray.scala 101:22]
  wire [2:0] _GEN_348 = _T_41 ? _GEN_331 : state; // @[Conditional.scala 39:67 PEArray.scala 100:22]
  wire [5:0] _GEN_353 = _T_31 ? _GEN_334 : _GEN_346; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_354 = _T_31 ? _GEN_330 : _GEN_347; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_355 = _T_31 ? _GEN_331 : _GEN_348; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_356 = _T_22 ? _GEN_330 : _GEN_354; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_357 = _T_22 ? _GEN_329 : _GEN_353; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_458 = _T_22 ? _GEN_331 : _GEN_355; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_690 = _T_3 ? _GEN_118 : {{2'd0}, GRU_out_width}; // @[Conditional.scala 40:58 PEArray.scala 104:26]
  FP16MulAdder FP16MAC ( // @[PEArray.scala 72:23]
    .io_a(FP16MAC_io_a),
    .io_b(FP16MAC_io_b),
    .io_c(FP16MAC_io_c),
    .io_out(FP16MAC_io_out)
  );
  assign io_ToRightPE = mux3out_reg; // @[PEArray.scala 95:16]
  assign io_ToBelowPE = mux2out_reg; // @[PEArray.scala 94:16]
  assign FP16MAC_io_a = sel1 ? io_FromL1 : io_FromLeftPE; // @[PEArray.scala 50:14 PEArray.scala 50:23 PEArray.scala 51:24]
  assign FP16MAC_io_b = sel5 ? mux4out : _GEN_105; // @[PEArray.scala 77:13 PEArray.scala 78:18 PEArray.scala 81:18]
  assign FP16MAC_io_c = sel5 ? _GEN_105 : mux4out; // @[PEArray.scala 77:13 PEArray.scala 79:18 PEArray.scala 82:18]
  always @(posedge clock) begin
    if (reset) begin // @[PEArray.scala 39:24]
      L0Index <= 6'h0; // @[PEArray.scala 39:24]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h2; // @[PEArray.scala 159:15]
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h4; // @[PEArray.scala 181:15]
      end else begin
        L0Index <= _GEN_357;
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_0 <= _GEN_229;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_1 <= _GEN_230;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_2 <= _GEN_231;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_3 <= _GEN_232;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_4 <= _GEN_233;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_5 <= _GEN_234;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_6 <= _GEN_235;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_7 <= _GEN_236;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_8 <= _GEN_237;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_9 <= _GEN_238;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_10 <= _GEN_239;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_11 <= _GEN_240;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_12 <= _GEN_241;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_13 <= _GEN_242;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_14 <= _GEN_243;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_15 <= _GEN_244;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_16 <= _GEN_245;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_17 <= _GEN_246;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_18 <= _GEN_247;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_19 <= _GEN_248;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_20 <= _GEN_249;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_21 <= _GEN_250;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_22 <= _GEN_251;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_23 <= _GEN_252;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_24 <= _GEN_253;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_25 <= _GEN_254;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_26 <= _GEN_255;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_27 <= _GEN_256;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_28 <= _GEN_257;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_29 <= _GEN_258;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_30 <= _GEN_259;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_31 <= _GEN_260;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_32 <= _GEN_261;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_33 <= _GEN_262;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_34 <= _GEN_263;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_35 <= _GEN_264;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_36 <= _GEN_265;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_37 <= _GEN_266;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_38 <= _GEN_267;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_39 <= _GEN_268;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_40 <= _GEN_269;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_41 <= _GEN_270;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_42 <= _GEN_271;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_43 <= _GEN_272;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_44 <= _GEN_273;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_45 <= _GEN_274;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_46 <= _GEN_275;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_47 <= _GEN_276;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_48 <= _GEN_277;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_49 <= _GEN_278;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_50 <= _GEN_279;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_51 <= _GEN_280;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_52 <= _GEN_281;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_53 <= _GEN_282;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_54 <= _GEN_283;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_55 <= _GEN_284;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_56 <= _GEN_285;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_57 <= _GEN_286;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_58 <= _GEN_287;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_59 <= _GEN_288;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_60 <= _GEN_289;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_61 <= _GEN_290;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_62 <= _GEN_291;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_63 <= _GEN_292;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_64 <= _GEN_293;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_65 <= _GEN_294;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_66 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_67 <= _GEN_296;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_68 <= _GEN_297;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_69 <= _GEN_298;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_70 <= _GEN_299;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_71 <= _GEN_300;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_72 <= _GEN_301;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_73 <= _GEN_302;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_74 <= _GEN_303;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_75 <= _GEN_304;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_76 <= _GEN_305;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_77 <= _GEN_306;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_78 <= _GEN_307;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_79 <= _GEN_308;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_80 <= _GEN_309;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_81 <= _GEN_310;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_82 <= _GEN_311;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_83 <= _GEN_312;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_84 <= _GEN_313;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_85 <= _GEN_314;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_86 <= _GEN_315;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_87 <= _GEN_316;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_88 <= _GEN_317;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_89 <= _GEN_318;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_90 <= _GEN_319;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_91 <= _GEN_320;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_92 <= _GEN_321;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_93 <= _GEN_322;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_94 <= _GEN_323;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_95 <= _GEN_324;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_96 <= _GEN_325;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_97 <= _GEN_326;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_98 <= _GEN_327;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_99 <= _GEN_328;
          end
        end
      end
    end
    if (reset) begin // @[PEArray.scala 100:22]
      state <= 3'h0; // @[PEArray.scala 100:22]
    end else if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[10]) begin // @[PEArray.scala 116:57]
        if (_T_6) begin // @[Conditional.scala 40:58]
          state <= 3'h0; // @[PEArray.scala 120:19]
        end else begin
          state <= _GEN_113;
        end
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      if (count == 10'h33) begin // @[PEArray.scala 164:27]
        state <= 3'h0; // @[PEArray.scala 166:15]
      end
    end else if (_T_16) begin // @[Conditional.scala 39:67]
      state <= _GEN_126;
    end else begin
      state <= _GEN_458;
    end
    if (reset) begin // @[PEArray.scala 90:28]
      mux2out_reg <= 16'h0; // @[PEArray.scala 90:28]
    end else begin
      mux2out_reg <= MAC_out; // @[PEArray.scala 90:28]
    end
    if (reset) begin // @[PEArray.scala 91:28]
      mux3out_reg <= 16'h0; // @[PEArray.scala 91:28]
    end else if (sel3) begin // @[PEArray.scala 56:14]
      mux3out_reg <= MAC_out; // @[PEArray.scala 56:23]
    end else if (sel1) begin // @[PEArray.scala 50:14]
      mux3out_reg <= io_FromL1; // @[PEArray.scala 50:23]
    end else begin
      mux3out_reg <= io_FromLeftPE; // @[PEArray.scala 51:24]
    end
    if (reset) begin // @[PEArray.scala 101:22]
      count <= 10'h0; // @[PEArray.scala 101:22]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        if (count == 10'h33) begin // @[PEArray.scala 164:27]
          count <= 10'h0; // @[PEArray.scala 165:15]
        end else begin
          count <= _GEN_120;
        end
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        count <= _GEN_125;
      end else begin
        count <= _GEN_356;
      end
    end
    if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[10]) begin // @[PEArray.scala 116:57]
        count_max <= io_control_signal_count; // @[PEArray.scala 143:19]
      end
    end
    if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[10]) begin // @[PEArray.scala 116:57]
        L0index_begin <= io_control_signal_L0index; // @[PEArray.scala 144:23]
      end
    end
    GRU_out_width <= _GEN_690[5:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  L0Index = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  L0Memory_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  L0Memory_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  L0Memory_2 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  L0Memory_3 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  L0Memory_4 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  L0Memory_5 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  L0Memory_6 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  L0Memory_7 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  L0Memory_8 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  L0Memory_9 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  L0Memory_10 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  L0Memory_11 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  L0Memory_12 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  L0Memory_13 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  L0Memory_14 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  L0Memory_15 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  L0Memory_16 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  L0Memory_17 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  L0Memory_18 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  L0Memory_19 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  L0Memory_20 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  L0Memory_21 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  L0Memory_22 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  L0Memory_23 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  L0Memory_24 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  L0Memory_25 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  L0Memory_26 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  L0Memory_27 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  L0Memory_28 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  L0Memory_29 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  L0Memory_30 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  L0Memory_31 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  L0Memory_32 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  L0Memory_33 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  L0Memory_34 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  L0Memory_35 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  L0Memory_36 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  L0Memory_37 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  L0Memory_38 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  L0Memory_39 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  L0Memory_40 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  L0Memory_41 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  L0Memory_42 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  L0Memory_43 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  L0Memory_44 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  L0Memory_45 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  L0Memory_46 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  L0Memory_47 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  L0Memory_48 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  L0Memory_49 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  L0Memory_50 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  L0Memory_51 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  L0Memory_52 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  L0Memory_53 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  L0Memory_54 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  L0Memory_55 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  L0Memory_56 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  L0Memory_57 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  L0Memory_58 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  L0Memory_59 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  L0Memory_60 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  L0Memory_61 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  L0Memory_62 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  L0Memory_63 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  L0Memory_64 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  L0Memory_65 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  L0Memory_66 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  L0Memory_67 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  L0Memory_68 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  L0Memory_69 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  L0Memory_70 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  L0Memory_71 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  L0Memory_72 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  L0Memory_73 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  L0Memory_74 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  L0Memory_75 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  L0Memory_76 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  L0Memory_77 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  L0Memory_78 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  L0Memory_79 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  L0Memory_80 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  L0Memory_81 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  L0Memory_82 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  L0Memory_83 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  L0Memory_84 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  L0Memory_85 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  L0Memory_86 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  L0Memory_87 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  L0Memory_88 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  L0Memory_89 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  L0Memory_90 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  L0Memory_91 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  L0Memory_92 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  L0Memory_93 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  L0Memory_94 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  L0Memory_95 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  L0Memory_96 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  L0Memory_97 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  L0Memory_98 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  L0Memory_99 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  state = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  mux2out_reg = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  mux3out_reg = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  count = _RAND_104[9:0];
  _RAND_105 = {1{`RANDOM}};
  count_max = _RAND_105[9:0];
  _RAND_106 = {1{`RANDOM}};
  L0index_begin = _RAND_106[5:0];
  _RAND_107 = {1{`RANDOM}};
  GRU_out_width = _RAND_107[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PE_6(
  input         clock,
  input         reset,
  input  [15:0] io_FromAbovePE,
  input  [15:0] io_FromLeftPE,
  input  [15:0] io_FromL1,
  input  [11:0] io_control_signal_mask,
  output [15:0] io_ToRightPE,
  output [15:0] io_ToBelowPE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] FP16MAC_io_a; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_b; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_c; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_out; // @[PEArray.scala 72:23]
  reg [5:0] L0Index; // @[PEArray.scala 39:24]
  reg [15:0] L0Memory_0; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_1; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_2; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_3; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_4; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_5; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_6; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_7; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_8; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_9; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_10; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_11; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_12; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_13; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_14; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_15; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_16; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_17; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_18; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_19; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_20; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_21; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_22; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_23; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_24; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_25; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_26; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_27; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_28; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_29; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_30; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_31; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_32; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_33; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_34; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_35; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_36; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_37; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_38; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_39; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_40; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_41; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_42; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_43; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_44; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_45; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_46; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_47; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_48; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_49; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_50; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_51; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_52; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_53; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_54; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_55; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_56; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_57; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_58; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_59; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_60; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_61; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_62; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_63; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_64; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_65; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_66; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_67; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_68; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_69; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_70; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_71; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_72; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_73; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_74; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_75; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_76; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_77; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_78; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_79; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_80; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_81; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_82; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_83; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_84; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_85; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_86; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_87; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_88; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_89; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_90; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_91; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_92; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_93; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_94; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_95; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_96; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_97; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_98; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_99; // @[PEArray.scala 40:21]
  reg [2:0] state; // @[PEArray.scala 100:22]
  wire  _T_3 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_12 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_16 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_22 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_31 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_41 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_342 = _T_41 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 231:12 PEArray.scala 32:8]
  wire  _GEN_349 = _T_31 ? 1'h0 : _GEN_342; // @[Conditional.scala 39:67 PEArray.scala 208:12]
  wire  _GEN_459 = _T_22 | _GEN_349; // @[Conditional.scala 39:67 PEArray.scala 32:8]
  wire  _GEN_463 = _T_16 ? 1'h0 : _GEN_459; // @[Conditional.scala 39:67]
  wire  _GEN_572 = _T_12 | _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 149:12]
  wire  sel1 = _T_3 | _GEN_572; // @[Conditional.scala 40:58 PEArray.scala 108:12]
  wire [15:0] MAC_out = FP16MAC_io_out; // @[PEArray.scala 47:21 PEArray.scala 85:11]
  wire  _GEN_465 = _T_16 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 177:12]
  wire  _GEN_580 = _T_12 | _GEN_465; // @[Conditional.scala 39:67 PEArray.scala 34:8]
  wire  sel3 = _T_3 | _GEN_580; // @[Conditional.scala 40:58 PEArray.scala 110:12]
  wire [1:0] _GEN_344 = _T_41 ? 2'h2 : 2'h0; // @[Conditional.scala 39:67 PEArray.scala 233:12 PEArray.scala 35:8]
  wire [1:0] _GEN_351 = _T_31 ? 2'h2 : _GEN_344; // @[Conditional.scala 39:67 PEArray.scala 210:12]
  wire [1:0] _GEN_461 = _T_22 ? 2'h0 : _GEN_351; // @[Conditional.scala 39:67 PEArray.scala 35:8]
  wire [1:0] _GEN_466 = _T_16 ? 2'h0 : _GEN_461; // @[Conditional.scala 39:67 PEArray.scala 178:12]
  wire [1:0] _GEN_574 = _T_12 ? 2'h0 : _GEN_466; // @[Conditional.scala 39:67]
  wire [1:0] sel4 = _T_3 ? 2'h0 : _GEN_574; // @[Conditional.scala 40:58 PEArray.scala 111:12]
  wire [15:0] _GEN_3 = sel4 == 2'h2 ? io_FromL1 : 16'h0; // @[PEArray.scala 65:28 PEArray.scala 66:15 PEArray.scala 69:15]
  wire [15:0] _GEN_4 = sel4 == 2'h1 ? io_FromAbovePE : _GEN_3; // @[PEArray.scala 62:28 PEArray.scala 63:15]
  wire [15:0] mux4out = sel4 == 2'h0 ? 16'h0 : _GEN_4; // @[PEArray.scala 59:22 PEArray.scala 60:13]
  wire [15:0] _GEN_7 = 6'h1 == L0Index ? L0Memory_1 : L0Memory_0; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_8 = 6'h2 == L0Index ? L0Memory_2 : _GEN_7; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_9 = 6'h3 == L0Index ? L0Memory_3 : _GEN_8; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_10 = 6'h4 == L0Index ? L0Memory_4 : _GEN_9; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_11 = 6'h5 == L0Index ? L0Memory_5 : _GEN_10; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_12 = 6'h6 == L0Index ? L0Memory_6 : _GEN_11; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_13 = 6'h7 == L0Index ? L0Memory_7 : _GEN_12; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_14 = 6'h8 == L0Index ? L0Memory_8 : _GEN_13; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_15 = 6'h9 == L0Index ? L0Memory_9 : _GEN_14; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_16 = 6'ha == L0Index ? L0Memory_10 : _GEN_15; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_17 = 6'hb == L0Index ? L0Memory_11 : _GEN_16; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_18 = 6'hc == L0Index ? L0Memory_12 : _GEN_17; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_19 = 6'hd == L0Index ? L0Memory_13 : _GEN_18; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_20 = 6'he == L0Index ? L0Memory_14 : _GEN_19; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_21 = 6'hf == L0Index ? L0Memory_15 : _GEN_20; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_22 = 6'h10 == L0Index ? L0Memory_16 : _GEN_21; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_23 = 6'h11 == L0Index ? L0Memory_17 : _GEN_22; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_24 = 6'h12 == L0Index ? L0Memory_18 : _GEN_23; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_25 = 6'h13 == L0Index ? L0Memory_19 : _GEN_24; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_26 = 6'h14 == L0Index ? L0Memory_20 : _GEN_25; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_27 = 6'h15 == L0Index ? L0Memory_21 : _GEN_26; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_28 = 6'h16 == L0Index ? L0Memory_22 : _GEN_27; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_29 = 6'h17 == L0Index ? L0Memory_23 : _GEN_28; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_30 = 6'h18 == L0Index ? L0Memory_24 : _GEN_29; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_31 = 6'h19 == L0Index ? L0Memory_25 : _GEN_30; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_32 = 6'h1a == L0Index ? L0Memory_26 : _GEN_31; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_33 = 6'h1b == L0Index ? L0Memory_27 : _GEN_32; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_34 = 6'h1c == L0Index ? L0Memory_28 : _GEN_33; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_35 = 6'h1d == L0Index ? L0Memory_29 : _GEN_34; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_36 = 6'h1e == L0Index ? L0Memory_30 : _GEN_35; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_37 = 6'h1f == L0Index ? L0Memory_31 : _GEN_36; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_38 = 6'h20 == L0Index ? L0Memory_32 : _GEN_37; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_39 = 6'h21 == L0Index ? L0Memory_33 : _GEN_38; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_40 = 6'h22 == L0Index ? L0Memory_34 : _GEN_39; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_41 = 6'h23 == L0Index ? L0Memory_35 : _GEN_40; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_42 = 6'h24 == L0Index ? L0Memory_36 : _GEN_41; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_43 = 6'h25 == L0Index ? L0Memory_37 : _GEN_42; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_44 = 6'h26 == L0Index ? L0Memory_38 : _GEN_43; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_45 = 6'h27 == L0Index ? L0Memory_39 : _GEN_44; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_46 = 6'h28 == L0Index ? L0Memory_40 : _GEN_45; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_47 = 6'h29 == L0Index ? L0Memory_41 : _GEN_46; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_48 = 6'h2a == L0Index ? L0Memory_42 : _GEN_47; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_49 = 6'h2b == L0Index ? L0Memory_43 : _GEN_48; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_50 = 6'h2c == L0Index ? L0Memory_44 : _GEN_49; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_51 = 6'h2d == L0Index ? L0Memory_45 : _GEN_50; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_52 = 6'h2e == L0Index ? L0Memory_46 : _GEN_51; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_53 = 6'h2f == L0Index ? L0Memory_47 : _GEN_52; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_54 = 6'h30 == L0Index ? L0Memory_48 : _GEN_53; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_55 = 6'h31 == L0Index ? L0Memory_49 : _GEN_54; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_56 = 6'h32 == L0Index ? L0Memory_50 : _GEN_55; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_57 = 6'h33 == L0Index ? L0Memory_51 : _GEN_56; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_58 = 6'h34 == L0Index ? L0Memory_52 : _GEN_57; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_59 = 6'h35 == L0Index ? L0Memory_53 : _GEN_58; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_60 = 6'h36 == L0Index ? L0Memory_54 : _GEN_59; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_61 = 6'h37 == L0Index ? L0Memory_55 : _GEN_60; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_62 = 6'h38 == L0Index ? L0Memory_56 : _GEN_61; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_63 = 6'h39 == L0Index ? L0Memory_57 : _GEN_62; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_64 = 6'h3a == L0Index ? L0Memory_58 : _GEN_63; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_65 = 6'h3b == L0Index ? L0Memory_59 : _GEN_64; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_66 = 6'h3c == L0Index ? L0Memory_60 : _GEN_65; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_67 = 6'h3d == L0Index ? L0Memory_61 : _GEN_66; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_68 = 6'h3e == L0Index ? L0Memory_62 : _GEN_67; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_69 = 6'h3f == L0Index ? L0Memory_63 : _GEN_68; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [6:0] _GEN_793 = {{1'd0}, L0Index}; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_70 = 7'h40 == _GEN_793 ? L0Memory_64 : _GEN_69; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_71 = 7'h41 == _GEN_793 ? L0Memory_65 : _GEN_70; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_72 = 7'h42 == _GEN_793 ? L0Memory_66 : _GEN_71; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_73 = 7'h43 == _GEN_793 ? L0Memory_67 : _GEN_72; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_74 = 7'h44 == _GEN_793 ? L0Memory_68 : _GEN_73; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_75 = 7'h45 == _GEN_793 ? L0Memory_69 : _GEN_74; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_76 = 7'h46 == _GEN_793 ? L0Memory_70 : _GEN_75; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_77 = 7'h47 == _GEN_793 ? L0Memory_71 : _GEN_76; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_78 = 7'h48 == _GEN_793 ? L0Memory_72 : _GEN_77; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_79 = 7'h49 == _GEN_793 ? L0Memory_73 : _GEN_78; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_80 = 7'h4a == _GEN_793 ? L0Memory_74 : _GEN_79; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_81 = 7'h4b == _GEN_793 ? L0Memory_75 : _GEN_80; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_82 = 7'h4c == _GEN_793 ? L0Memory_76 : _GEN_81; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_83 = 7'h4d == _GEN_793 ? L0Memory_77 : _GEN_82; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_84 = 7'h4e == _GEN_793 ? L0Memory_78 : _GEN_83; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_85 = 7'h4f == _GEN_793 ? L0Memory_79 : _GEN_84; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_86 = 7'h50 == _GEN_793 ? L0Memory_80 : _GEN_85; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_87 = 7'h51 == _GEN_793 ? L0Memory_81 : _GEN_86; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_88 = 7'h52 == _GEN_793 ? L0Memory_82 : _GEN_87; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_89 = 7'h53 == _GEN_793 ? L0Memory_83 : _GEN_88; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_90 = 7'h54 == _GEN_793 ? L0Memory_84 : _GEN_89; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_91 = 7'h55 == _GEN_793 ? L0Memory_85 : _GEN_90; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_92 = 7'h56 == _GEN_793 ? L0Memory_86 : _GEN_91; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_93 = 7'h57 == _GEN_793 ? L0Memory_87 : _GEN_92; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_94 = 7'h58 == _GEN_793 ? L0Memory_88 : _GEN_93; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_95 = 7'h59 == _GEN_793 ? L0Memory_89 : _GEN_94; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_96 = 7'h5a == _GEN_793 ? L0Memory_90 : _GEN_95; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_97 = 7'h5b == _GEN_793 ? L0Memory_91 : _GEN_96; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_98 = 7'h5c == _GEN_793 ? L0Memory_92 : _GEN_97; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_99 = 7'h5d == _GEN_793 ? L0Memory_93 : _GEN_98; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_100 = 7'h5e == _GEN_793 ? L0Memory_94 : _GEN_99; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_101 = 7'h5f == _GEN_793 ? L0Memory_95 : _GEN_100; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_102 = 7'h60 == _GEN_793 ? L0Memory_96 : _GEN_101; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_103 = 7'h61 == _GEN_793 ? L0Memory_97 : _GEN_102; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_104 = 7'h62 == _GEN_793 ? L0Memory_98 : _GEN_103; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_105 = 7'h63 == _GEN_793 ? L0Memory_99 : _GEN_104; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire  _GEN_575 = _T_12 ? 1'h0 : _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 157:12]
  wire  sel5 = _T_3 ? 1'h0 : _GEN_575; // @[Conditional.scala 40:58 PEArray.scala 112:12]
  reg [15:0] mux2out_reg; // @[PEArray.scala 90:28]
  reg [15:0] mux3out_reg; // @[PEArray.scala 91:28]
  reg [9:0] count; // @[PEArray.scala 101:22]
  reg [5:0] GRU_out_width; // @[PEArray.scala 104:26]
  wire [7:0] _GEN_118 = io_control_signal_mask[9] ? 8'h0 : {{2'd0}, GRU_out_width}; // @[PEArray.scala 116:57 PEArray.scala 145:23 PEArray.scala 104:26]
  wire [9:0] _count_T_1 = count + 10'h1; // @[PEArray.scala 162:24]
  wire [9:0] _GEN_120 = count != 10'h33 ? _count_T_1 : count; // @[PEArray.scala 161:27 PEArray.scala 162:15 PEArray.scala 101:22]
  wire [9:0] _GEN_124 = count != 10'h188 ? _count_T_1 : count; // @[PEArray.scala 183:28 PEArray.scala 184:15 PEArray.scala 101:22]
  wire [9:0] _GEN_125 = count == 10'h188 ? 10'h0 : _GEN_124; // @[PEArray.scala 186:28 PEArray.scala 187:15]
  wire [2:0] _GEN_126 = count == 10'h188 ? 3'h0 : state; // @[PEArray.scala 186:28 PEArray.scala 188:15 PEArray.scala 100:22]
  wire [9:0] _GEN_127 = count != 10'h0 ? _count_T_1 : count; // @[PEArray.scala 192:32 PEArray.scala 193:15 PEArray.scala 101:22]
  wire  _T_24 = count == 10'h0; // @[PEArray.scala 195:18]
  wire [5:0] _GEN_128 = count == 10'h0 ? 6'h0 : L0Index; // @[PEArray.scala 195:26 PEArray.scala 196:17 PEArray.scala 39:24]
  wire [9:0] _T_27 = 10'h0 - 10'h1; // @[PEArray.scala 198:51]
  wire [15:0] _GEN_129 = 6'h0 == L0Index ? io_FromL1 : L0Memory_0; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_130 = 6'h1 == L0Index ? io_FromL1 : L0Memory_1; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_131 = 6'h2 == L0Index ? io_FromL1 : L0Memory_2; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_132 = 6'h3 == L0Index ? io_FromL1 : L0Memory_3; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_133 = 6'h4 == L0Index ? io_FromL1 : L0Memory_4; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_134 = 6'h5 == L0Index ? io_FromL1 : L0Memory_5; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_135 = 6'h6 == L0Index ? io_FromL1 : L0Memory_6; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_136 = 6'h7 == L0Index ? io_FromL1 : L0Memory_7; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_137 = 6'h8 == L0Index ? io_FromL1 : L0Memory_8; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_138 = 6'h9 == L0Index ? io_FromL1 : L0Memory_9; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_139 = 6'ha == L0Index ? io_FromL1 : L0Memory_10; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_140 = 6'hb == L0Index ? io_FromL1 : L0Memory_11; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_141 = 6'hc == L0Index ? io_FromL1 : L0Memory_12; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_142 = 6'hd == L0Index ? io_FromL1 : L0Memory_13; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_143 = 6'he == L0Index ? io_FromL1 : L0Memory_14; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_144 = 6'hf == L0Index ? io_FromL1 : L0Memory_15; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_145 = 6'h10 == L0Index ? io_FromL1 : L0Memory_16; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_146 = 6'h11 == L0Index ? io_FromL1 : L0Memory_17; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_147 = 6'h12 == L0Index ? io_FromL1 : L0Memory_18; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_148 = 6'h13 == L0Index ? io_FromL1 : L0Memory_19; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_149 = 6'h14 == L0Index ? io_FromL1 : L0Memory_20; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_150 = 6'h15 == L0Index ? io_FromL1 : L0Memory_21; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_151 = 6'h16 == L0Index ? io_FromL1 : L0Memory_22; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_152 = 6'h17 == L0Index ? io_FromL1 : L0Memory_23; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_153 = 6'h18 == L0Index ? io_FromL1 : L0Memory_24; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_154 = 6'h19 == L0Index ? io_FromL1 : L0Memory_25; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_155 = 6'h1a == L0Index ? io_FromL1 : L0Memory_26; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_156 = 6'h1b == L0Index ? io_FromL1 : L0Memory_27; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_157 = 6'h1c == L0Index ? io_FromL1 : L0Memory_28; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_158 = 6'h1d == L0Index ? io_FromL1 : L0Memory_29; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_159 = 6'h1e == L0Index ? io_FromL1 : L0Memory_30; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_160 = 6'h1f == L0Index ? io_FromL1 : L0Memory_31; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_161 = 6'h20 == L0Index ? io_FromL1 : L0Memory_32; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_162 = 6'h21 == L0Index ? io_FromL1 : L0Memory_33; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_163 = 6'h22 == L0Index ? io_FromL1 : L0Memory_34; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_164 = 6'h23 == L0Index ? io_FromL1 : L0Memory_35; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_165 = 6'h24 == L0Index ? io_FromL1 : L0Memory_36; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_166 = 6'h25 == L0Index ? io_FromL1 : L0Memory_37; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_167 = 6'h26 == L0Index ? io_FromL1 : L0Memory_38; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_168 = 6'h27 == L0Index ? io_FromL1 : L0Memory_39; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_169 = 6'h28 == L0Index ? io_FromL1 : L0Memory_40; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_170 = 6'h29 == L0Index ? io_FromL1 : L0Memory_41; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_171 = 6'h2a == L0Index ? io_FromL1 : L0Memory_42; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_172 = 6'h2b == L0Index ? io_FromL1 : L0Memory_43; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_173 = 6'h2c == L0Index ? io_FromL1 : L0Memory_44; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_174 = 6'h2d == L0Index ? io_FromL1 : L0Memory_45; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_175 = 6'h2e == L0Index ? io_FromL1 : L0Memory_46; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_176 = 6'h2f == L0Index ? io_FromL1 : L0Memory_47; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_177 = 6'h30 == L0Index ? io_FromL1 : L0Memory_48; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_178 = 6'h31 == L0Index ? io_FromL1 : L0Memory_49; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_179 = 6'h32 == L0Index ? io_FromL1 : L0Memory_50; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_180 = 6'h33 == L0Index ? io_FromL1 : L0Memory_51; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_181 = 6'h34 == L0Index ? io_FromL1 : L0Memory_52; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_182 = 6'h35 == L0Index ? io_FromL1 : L0Memory_53; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_183 = 6'h36 == L0Index ? io_FromL1 : L0Memory_54; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_184 = 6'h37 == L0Index ? io_FromL1 : L0Memory_55; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_185 = 6'h38 == L0Index ? io_FromL1 : L0Memory_56; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_186 = 6'h39 == L0Index ? io_FromL1 : L0Memory_57; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_187 = 6'h3a == L0Index ? io_FromL1 : L0Memory_58; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_188 = 6'h3b == L0Index ? io_FromL1 : L0Memory_59; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_189 = 6'h3c == L0Index ? io_FromL1 : L0Memory_60; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_190 = 6'h3d == L0Index ? io_FromL1 : L0Memory_61; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_191 = 6'h3e == L0Index ? io_FromL1 : L0Memory_62; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_192 = 6'h3f == L0Index ? io_FromL1 : L0Memory_63; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_193 = 7'h40 == _GEN_793 ? io_FromL1 : L0Memory_64; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_194 = 7'h41 == _GEN_793 ? io_FromL1 : L0Memory_65; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_195 = 7'h42 == _GEN_793 ? io_FromL1 : L0Memory_66; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_196 = 7'h43 == _GEN_793 ? io_FromL1 : L0Memory_67; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_197 = 7'h44 == _GEN_793 ? io_FromL1 : L0Memory_68; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_198 = 7'h45 == _GEN_793 ? io_FromL1 : L0Memory_69; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_199 = 7'h46 == _GEN_793 ? io_FromL1 : L0Memory_70; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_200 = 7'h47 == _GEN_793 ? io_FromL1 : L0Memory_71; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_201 = 7'h48 == _GEN_793 ? io_FromL1 : L0Memory_72; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_202 = 7'h49 == _GEN_793 ? io_FromL1 : L0Memory_73; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_203 = 7'h4a == _GEN_793 ? io_FromL1 : L0Memory_74; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_204 = 7'h4b == _GEN_793 ? io_FromL1 : L0Memory_75; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_205 = 7'h4c == _GEN_793 ? io_FromL1 : L0Memory_76; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_206 = 7'h4d == _GEN_793 ? io_FromL1 : L0Memory_77; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_207 = 7'h4e == _GEN_793 ? io_FromL1 : L0Memory_78; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_208 = 7'h4f == _GEN_793 ? io_FromL1 : L0Memory_79; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_209 = 7'h50 == _GEN_793 ? io_FromL1 : L0Memory_80; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_210 = 7'h51 == _GEN_793 ? io_FromL1 : L0Memory_81; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_211 = 7'h52 == _GEN_793 ? io_FromL1 : L0Memory_82; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_212 = 7'h53 == _GEN_793 ? io_FromL1 : L0Memory_83; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_213 = 7'h54 == _GEN_793 ? io_FromL1 : L0Memory_84; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_214 = 7'h55 == _GEN_793 ? io_FromL1 : L0Memory_85; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_215 = 7'h56 == _GEN_793 ? io_FromL1 : L0Memory_86; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_216 = 7'h57 == _GEN_793 ? io_FromL1 : L0Memory_87; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_217 = 7'h58 == _GEN_793 ? io_FromL1 : L0Memory_88; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_218 = 7'h59 == _GEN_793 ? io_FromL1 : L0Memory_89; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_219 = 7'h5a == _GEN_793 ? io_FromL1 : L0Memory_90; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_220 = 7'h5b == _GEN_793 ? io_FromL1 : L0Memory_91; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_221 = 7'h5c == _GEN_793 ? io_FromL1 : L0Memory_92; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_222 = 7'h5d == _GEN_793 ? io_FromL1 : L0Memory_93; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_223 = 7'h5e == _GEN_793 ? io_FromL1 : L0Memory_94; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_224 = 7'h5f == _GEN_793 ? io_FromL1 : L0Memory_95; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_225 = 7'h60 == _GEN_793 ? io_FromL1 : L0Memory_96; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_226 = 7'h61 == _GEN_793 ? io_FromL1 : L0Memory_97; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_227 = 7'h62 == _GEN_793 ? io_FromL1 : L0Memory_98; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_228 = 7'h63 == _GEN_793 ? io_FromL1 : L0Memory_99; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [5:0] _L0Index_T_2 = L0Index + 6'h1; // @[PEArray.scala 200:28]
  wire [15:0] _GEN_229 = count >= 10'h1 & count <= _T_27 ? _GEN_129 : L0Memory_0; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_230 = count >= 10'h1 & count <= _T_27 ? _GEN_130 : L0Memory_1; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_231 = count >= 10'h1 & count <= _T_27 ? _GEN_131 : L0Memory_2; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_232 = count >= 10'h1 & count <= _T_27 ? _GEN_132 : L0Memory_3; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_233 = count >= 10'h1 & count <= _T_27 ? _GEN_133 : L0Memory_4; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_234 = count >= 10'h1 & count <= _T_27 ? _GEN_134 : L0Memory_5; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_235 = count >= 10'h1 & count <= _T_27 ? _GEN_135 : L0Memory_6; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_236 = count >= 10'h1 & count <= _T_27 ? _GEN_136 : L0Memory_7; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_237 = count >= 10'h1 & count <= _T_27 ? _GEN_137 : L0Memory_8; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_238 = count >= 10'h1 & count <= _T_27 ? _GEN_138 : L0Memory_9; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_239 = count >= 10'h1 & count <= _T_27 ? _GEN_139 : L0Memory_10; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_240 = count >= 10'h1 & count <= _T_27 ? _GEN_140 : L0Memory_11; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_241 = count >= 10'h1 & count <= _T_27 ? _GEN_141 : L0Memory_12; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_242 = count >= 10'h1 & count <= _T_27 ? _GEN_142 : L0Memory_13; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_243 = count >= 10'h1 & count <= _T_27 ? _GEN_143 : L0Memory_14; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_244 = count >= 10'h1 & count <= _T_27 ? _GEN_144 : L0Memory_15; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_245 = count >= 10'h1 & count <= _T_27 ? _GEN_145 : L0Memory_16; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_246 = count >= 10'h1 & count <= _T_27 ? _GEN_146 : L0Memory_17; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_247 = count >= 10'h1 & count <= _T_27 ? _GEN_147 : L0Memory_18; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_248 = count >= 10'h1 & count <= _T_27 ? _GEN_148 : L0Memory_19; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_249 = count >= 10'h1 & count <= _T_27 ? _GEN_149 : L0Memory_20; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_250 = count >= 10'h1 & count <= _T_27 ? _GEN_150 : L0Memory_21; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_251 = count >= 10'h1 & count <= _T_27 ? _GEN_151 : L0Memory_22; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_252 = count >= 10'h1 & count <= _T_27 ? _GEN_152 : L0Memory_23; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_253 = count >= 10'h1 & count <= _T_27 ? _GEN_153 : L0Memory_24; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_254 = count >= 10'h1 & count <= _T_27 ? _GEN_154 : L0Memory_25; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_255 = count >= 10'h1 & count <= _T_27 ? _GEN_155 : L0Memory_26; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_256 = count >= 10'h1 & count <= _T_27 ? _GEN_156 : L0Memory_27; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_257 = count >= 10'h1 & count <= _T_27 ? _GEN_157 : L0Memory_28; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_258 = count >= 10'h1 & count <= _T_27 ? _GEN_158 : L0Memory_29; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_259 = count >= 10'h1 & count <= _T_27 ? _GEN_159 : L0Memory_30; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_260 = count >= 10'h1 & count <= _T_27 ? _GEN_160 : L0Memory_31; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_261 = count >= 10'h1 & count <= _T_27 ? _GEN_161 : L0Memory_32; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_262 = count >= 10'h1 & count <= _T_27 ? _GEN_162 : L0Memory_33; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_263 = count >= 10'h1 & count <= _T_27 ? _GEN_163 : L0Memory_34; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_264 = count >= 10'h1 & count <= _T_27 ? _GEN_164 : L0Memory_35; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_265 = count >= 10'h1 & count <= _T_27 ? _GEN_165 : L0Memory_36; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_266 = count >= 10'h1 & count <= _T_27 ? _GEN_166 : L0Memory_37; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_267 = count >= 10'h1 & count <= _T_27 ? _GEN_167 : L0Memory_38; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_268 = count >= 10'h1 & count <= _T_27 ? _GEN_168 : L0Memory_39; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_269 = count >= 10'h1 & count <= _T_27 ? _GEN_169 : L0Memory_40; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_270 = count >= 10'h1 & count <= _T_27 ? _GEN_170 : L0Memory_41; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_271 = count >= 10'h1 & count <= _T_27 ? _GEN_171 : L0Memory_42; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_272 = count >= 10'h1 & count <= _T_27 ? _GEN_172 : L0Memory_43; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_273 = count >= 10'h1 & count <= _T_27 ? _GEN_173 : L0Memory_44; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_274 = count >= 10'h1 & count <= _T_27 ? _GEN_174 : L0Memory_45; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_275 = count >= 10'h1 & count <= _T_27 ? _GEN_175 : L0Memory_46; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_276 = count >= 10'h1 & count <= _T_27 ? _GEN_176 : L0Memory_47; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_277 = count >= 10'h1 & count <= _T_27 ? _GEN_177 : L0Memory_48; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_278 = count >= 10'h1 & count <= _T_27 ? _GEN_178 : L0Memory_49; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_279 = count >= 10'h1 & count <= _T_27 ? _GEN_179 : L0Memory_50; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_280 = count >= 10'h1 & count <= _T_27 ? _GEN_180 : L0Memory_51; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_281 = count >= 10'h1 & count <= _T_27 ? _GEN_181 : L0Memory_52; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_282 = count >= 10'h1 & count <= _T_27 ? _GEN_182 : L0Memory_53; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_283 = count >= 10'h1 & count <= _T_27 ? _GEN_183 : L0Memory_54; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_284 = count >= 10'h1 & count <= _T_27 ? _GEN_184 : L0Memory_55; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_285 = count >= 10'h1 & count <= _T_27 ? _GEN_185 : L0Memory_56; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_286 = count >= 10'h1 & count <= _T_27 ? _GEN_186 : L0Memory_57; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_287 = count >= 10'h1 & count <= _T_27 ? _GEN_187 : L0Memory_58; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_288 = count >= 10'h1 & count <= _T_27 ? _GEN_188 : L0Memory_59; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_289 = count >= 10'h1 & count <= _T_27 ? _GEN_189 : L0Memory_60; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_290 = count >= 10'h1 & count <= _T_27 ? _GEN_190 : L0Memory_61; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_291 = count >= 10'h1 & count <= _T_27 ? _GEN_191 : L0Memory_62; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_292 = count >= 10'h1 & count <= _T_27 ? _GEN_192 : L0Memory_63; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_293 = count >= 10'h1 & count <= _T_27 ? _GEN_193 : L0Memory_64; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_294 = count >= 10'h1 & count <= _T_27 ? _GEN_194 : L0Memory_65; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_295 = count >= 10'h1 & count <= _T_27 ? _GEN_195 : L0Memory_66; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_296 = count >= 10'h1 & count <= _T_27 ? _GEN_196 : L0Memory_67; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_297 = count >= 10'h1 & count <= _T_27 ? _GEN_197 : L0Memory_68; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_298 = count >= 10'h1 & count <= _T_27 ? _GEN_198 : L0Memory_69; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_299 = count >= 10'h1 & count <= _T_27 ? _GEN_199 : L0Memory_70; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_300 = count >= 10'h1 & count <= _T_27 ? _GEN_200 : L0Memory_71; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_301 = count >= 10'h1 & count <= _T_27 ? _GEN_201 : L0Memory_72; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_302 = count >= 10'h1 & count <= _T_27 ? _GEN_202 : L0Memory_73; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_303 = count >= 10'h1 & count <= _T_27 ? _GEN_203 : L0Memory_74; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_304 = count >= 10'h1 & count <= _T_27 ? _GEN_204 : L0Memory_75; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_305 = count >= 10'h1 & count <= _T_27 ? _GEN_205 : L0Memory_76; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_306 = count >= 10'h1 & count <= _T_27 ? _GEN_206 : L0Memory_77; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_307 = count >= 10'h1 & count <= _T_27 ? _GEN_207 : L0Memory_78; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_308 = count >= 10'h1 & count <= _T_27 ? _GEN_208 : L0Memory_79; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_309 = count >= 10'h1 & count <= _T_27 ? _GEN_209 : L0Memory_80; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_310 = count >= 10'h1 & count <= _T_27 ? _GEN_210 : L0Memory_81; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_311 = count >= 10'h1 & count <= _T_27 ? _GEN_211 : L0Memory_82; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_312 = count >= 10'h1 & count <= _T_27 ? _GEN_212 : L0Memory_83; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_313 = count >= 10'h1 & count <= _T_27 ? _GEN_213 : L0Memory_84; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_314 = count >= 10'h1 & count <= _T_27 ? _GEN_214 : L0Memory_85; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_315 = count >= 10'h1 & count <= _T_27 ? _GEN_215 : L0Memory_86; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_316 = count >= 10'h1 & count <= _T_27 ? _GEN_216 : L0Memory_87; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_317 = count >= 10'h1 & count <= _T_27 ? _GEN_217 : L0Memory_88; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_318 = count >= 10'h1 & count <= _T_27 ? _GEN_218 : L0Memory_89; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_319 = count >= 10'h1 & count <= _T_27 ? _GEN_219 : L0Memory_90; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_320 = count >= 10'h1 & count <= _T_27 ? _GEN_220 : L0Memory_91; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_321 = count >= 10'h1 & count <= _T_27 ? _GEN_221 : L0Memory_92; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_322 = count >= 10'h1 & count <= _T_27 ? _GEN_222 : L0Memory_93; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_323 = count >= 10'h1 & count <= _T_27 ? _GEN_223 : L0Memory_94; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_324 = count >= 10'h1 & count <= _T_27 ? _GEN_224 : L0Memory_95; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_325 = count >= 10'h1 & count <= _T_27 ? _GEN_225 : L0Memory_96; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_326 = count >= 10'h1 & count <= _T_27 ? _GEN_226 : L0Memory_97; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_327 = count >= 10'h1 & count <= _T_27 ? _GEN_227 : L0Memory_98; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_328 = count >= 10'h1 & count <= _T_27 ? _GEN_228 : L0Memory_99; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [5:0] _GEN_329 = count >= 10'h1 & count <= _T_27 ? _L0Index_T_2 : _GEN_128; // @[PEArray.scala 198:59 PEArray.scala 200:17]
  wire [9:0] _GEN_330 = _T_24 ? 10'h0 : _GEN_127; // @[PEArray.scala 202:32 PEArray.scala 203:15]
  wire [2:0] _GEN_331 = _T_24 ? 3'h0 : state; // @[PEArray.scala 202:32 PEArray.scala 204:15 PEArray.scala 100:22]
  wire [9:0] _GEN_865 = {{4'd0}, GRU_out_width}; // @[PEArray.scala 220:19]
  wire [9:0] _GEN_0 = count % _GEN_865; // @[PEArray.scala 220:19]
  wire [5:0] _T_36 = _GEN_0[5:0]; // @[PEArray.scala 220:19]
  wire [5:0] _T_38 = GRU_out_width - 6'h1; // @[PEArray.scala 220:55]
  wire [5:0] _GEN_334 = _T_36 == _T_38 ? _L0Index_T_2 : 6'h0; // @[PEArray.scala 220:62 PEArray.scala 221:17 PEArray.scala 214:15]
  wire [5:0] _GEN_346 = _T_41 ? _GEN_334 : L0Index; // @[Conditional.scala 39:67 PEArray.scala 39:24]
  wire [9:0] _GEN_347 = _T_41 ? _GEN_330 : count; // @[Conditional.scala 39:67 PEArray.scala 101:22]
  wire [2:0] _GEN_348 = _T_41 ? _GEN_331 : state; // @[Conditional.scala 39:67 PEArray.scala 100:22]
  wire [5:0] _GEN_353 = _T_31 ? _GEN_334 : _GEN_346; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_354 = _T_31 ? _GEN_330 : _GEN_347; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_355 = _T_31 ? _GEN_331 : _GEN_348; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_356 = _T_22 ? _GEN_330 : _GEN_354; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_357 = _T_22 ? _GEN_329 : _GEN_353; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_458 = _T_22 ? _GEN_331 : _GEN_355; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_690 = _T_3 ? _GEN_118 : {{2'd0}, GRU_out_width}; // @[Conditional.scala 40:58 PEArray.scala 104:26]
  FP16MulAdder FP16MAC ( // @[PEArray.scala 72:23]
    .io_a(FP16MAC_io_a),
    .io_b(FP16MAC_io_b),
    .io_c(FP16MAC_io_c),
    .io_out(FP16MAC_io_out)
  );
  assign io_ToRightPE = mux3out_reg; // @[PEArray.scala 95:16]
  assign io_ToBelowPE = mux2out_reg; // @[PEArray.scala 94:16]
  assign FP16MAC_io_a = sel1 ? io_FromL1 : io_FromLeftPE; // @[PEArray.scala 50:14 PEArray.scala 50:23 PEArray.scala 51:24]
  assign FP16MAC_io_b = sel5 ? mux4out : _GEN_105; // @[PEArray.scala 77:13 PEArray.scala 78:18 PEArray.scala 81:18]
  assign FP16MAC_io_c = sel5 ? _GEN_105 : mux4out; // @[PEArray.scala 77:13 PEArray.scala 79:18 PEArray.scala 82:18]
  always @(posedge clock) begin
    if (reset) begin // @[PEArray.scala 39:24]
      L0Index <= 6'h0; // @[PEArray.scala 39:24]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h0; // @[PEArray.scala 159:15]
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h5; // @[PEArray.scala 181:15]
      end else begin
        L0Index <= _GEN_357;
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_0 <= _GEN_229;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_1 <= _GEN_230;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_2 <= _GEN_231;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_3 <= _GEN_232;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_4 <= _GEN_233;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_5 <= _GEN_234;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_6 <= _GEN_235;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_7 <= _GEN_236;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_8 <= _GEN_237;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_9 <= _GEN_238;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_10 <= _GEN_239;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_11 <= _GEN_240;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_12 <= _GEN_241;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_13 <= _GEN_242;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_14 <= _GEN_243;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_15 <= _GEN_244;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_16 <= _GEN_245;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_17 <= _GEN_246;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_18 <= _GEN_247;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_19 <= _GEN_248;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_20 <= _GEN_249;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_21 <= _GEN_250;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_22 <= _GEN_251;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_23 <= _GEN_252;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_24 <= _GEN_253;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_25 <= _GEN_254;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_26 <= _GEN_255;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_27 <= _GEN_256;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_28 <= _GEN_257;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_29 <= _GEN_258;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_30 <= _GEN_259;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_31 <= _GEN_260;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_32 <= _GEN_261;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_33 <= _GEN_262;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_34 <= _GEN_263;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_35 <= _GEN_264;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_36 <= _GEN_265;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_37 <= _GEN_266;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_38 <= _GEN_267;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_39 <= _GEN_268;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_40 <= _GEN_269;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_41 <= _GEN_270;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_42 <= _GEN_271;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_43 <= _GEN_272;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_44 <= _GEN_273;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_45 <= _GEN_274;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_46 <= _GEN_275;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_47 <= _GEN_276;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_48 <= _GEN_277;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_49 <= _GEN_278;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_50 <= _GEN_279;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_51 <= _GEN_280;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_52 <= _GEN_281;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_53 <= _GEN_282;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_54 <= _GEN_283;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_55 <= _GEN_284;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_56 <= _GEN_285;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_57 <= _GEN_286;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_58 <= _GEN_287;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_59 <= _GEN_288;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_60 <= _GEN_289;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_61 <= _GEN_290;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_62 <= _GEN_291;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_63 <= _GEN_292;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_64 <= _GEN_293;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_65 <= _GEN_294;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_66 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_67 <= _GEN_296;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_68 <= _GEN_297;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_69 <= _GEN_298;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_70 <= _GEN_299;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_71 <= _GEN_300;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_72 <= _GEN_301;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_73 <= _GEN_302;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_74 <= _GEN_303;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_75 <= _GEN_304;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_76 <= _GEN_305;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_77 <= _GEN_306;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_78 <= _GEN_307;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_79 <= _GEN_308;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_80 <= _GEN_309;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_81 <= _GEN_310;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_82 <= _GEN_311;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_83 <= _GEN_312;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_84 <= _GEN_313;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_85 <= _GEN_314;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_86 <= _GEN_315;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_87 <= _GEN_316;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_88 <= _GEN_317;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_89 <= _GEN_318;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_90 <= _GEN_319;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_91 <= _GEN_320;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_92 <= _GEN_321;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_93 <= _GEN_322;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_94 <= _GEN_323;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_95 <= _GEN_324;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_96 <= _GEN_325;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_97 <= _GEN_326;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_98 <= _GEN_327;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_99 <= _GEN_328;
          end
        end
      end
    end
    if (reset) begin // @[PEArray.scala 100:22]
      state <= 3'h0; // @[PEArray.scala 100:22]
    end else if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[9]) begin // @[PEArray.scala 116:57]
        state <= 3'h1;
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      if (count == 10'h33) begin // @[PEArray.scala 164:27]
        state <= 3'h0; // @[PEArray.scala 166:15]
      end
    end else if (_T_16) begin // @[Conditional.scala 39:67]
      state <= _GEN_126;
    end else begin
      state <= _GEN_458;
    end
    if (reset) begin // @[PEArray.scala 90:28]
      mux2out_reg <= 16'h0; // @[PEArray.scala 90:28]
    end else begin
      mux2out_reg <= MAC_out; // @[PEArray.scala 90:28]
    end
    if (reset) begin // @[PEArray.scala 91:28]
      mux3out_reg <= 16'h0; // @[PEArray.scala 91:28]
    end else if (sel3) begin // @[PEArray.scala 56:14]
      mux3out_reg <= MAC_out; // @[PEArray.scala 56:23]
    end else if (sel1) begin // @[PEArray.scala 50:14]
      mux3out_reg <= io_FromL1; // @[PEArray.scala 50:23]
    end else begin
      mux3out_reg <= io_FromLeftPE; // @[PEArray.scala 51:24]
    end
    if (reset) begin // @[PEArray.scala 101:22]
      count <= 10'h0; // @[PEArray.scala 101:22]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        if (count == 10'h33) begin // @[PEArray.scala 164:27]
          count <= 10'h0; // @[PEArray.scala 165:15]
        end else begin
          count <= _GEN_120;
        end
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        count <= _GEN_125;
      end else begin
        count <= _GEN_356;
      end
    end
    GRU_out_width <= _GEN_690[5:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  L0Index = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  L0Memory_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  L0Memory_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  L0Memory_2 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  L0Memory_3 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  L0Memory_4 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  L0Memory_5 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  L0Memory_6 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  L0Memory_7 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  L0Memory_8 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  L0Memory_9 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  L0Memory_10 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  L0Memory_11 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  L0Memory_12 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  L0Memory_13 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  L0Memory_14 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  L0Memory_15 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  L0Memory_16 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  L0Memory_17 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  L0Memory_18 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  L0Memory_19 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  L0Memory_20 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  L0Memory_21 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  L0Memory_22 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  L0Memory_23 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  L0Memory_24 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  L0Memory_25 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  L0Memory_26 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  L0Memory_27 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  L0Memory_28 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  L0Memory_29 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  L0Memory_30 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  L0Memory_31 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  L0Memory_32 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  L0Memory_33 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  L0Memory_34 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  L0Memory_35 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  L0Memory_36 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  L0Memory_37 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  L0Memory_38 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  L0Memory_39 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  L0Memory_40 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  L0Memory_41 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  L0Memory_42 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  L0Memory_43 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  L0Memory_44 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  L0Memory_45 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  L0Memory_46 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  L0Memory_47 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  L0Memory_48 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  L0Memory_49 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  L0Memory_50 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  L0Memory_51 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  L0Memory_52 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  L0Memory_53 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  L0Memory_54 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  L0Memory_55 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  L0Memory_56 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  L0Memory_57 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  L0Memory_58 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  L0Memory_59 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  L0Memory_60 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  L0Memory_61 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  L0Memory_62 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  L0Memory_63 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  L0Memory_64 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  L0Memory_65 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  L0Memory_66 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  L0Memory_67 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  L0Memory_68 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  L0Memory_69 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  L0Memory_70 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  L0Memory_71 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  L0Memory_72 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  L0Memory_73 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  L0Memory_74 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  L0Memory_75 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  L0Memory_76 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  L0Memory_77 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  L0Memory_78 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  L0Memory_79 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  L0Memory_80 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  L0Memory_81 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  L0Memory_82 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  L0Memory_83 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  L0Memory_84 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  L0Memory_85 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  L0Memory_86 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  L0Memory_87 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  L0Memory_88 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  L0Memory_89 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  L0Memory_90 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  L0Memory_91 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  L0Memory_92 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  L0Memory_93 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  L0Memory_94 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  L0Memory_95 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  L0Memory_96 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  L0Memory_97 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  L0Memory_98 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  L0Memory_99 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  state = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  mux2out_reg = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  mux3out_reg = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  count = _RAND_104[9:0];
  _RAND_105 = {1{`RANDOM}};
  GRU_out_width = _RAND_105[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PE_7(
  input         clock,
  input         reset,
  input  [15:0] io_FromAbovePE,
  input  [15:0] io_FromLeftPE,
  input  [15:0] io_FromL1,
  input  [11:0] io_control_signal_mask,
  output [15:0] io_ToRightPE,
  output [15:0] io_ToBelowPE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] FP16MAC_io_a; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_b; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_c; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_out; // @[PEArray.scala 72:23]
  reg [5:0] L0Index; // @[PEArray.scala 39:24]
  reg [15:0] L0Memory_0; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_1; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_2; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_3; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_4; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_5; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_6; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_7; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_8; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_9; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_10; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_11; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_12; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_13; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_14; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_15; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_16; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_17; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_18; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_19; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_20; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_21; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_22; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_23; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_24; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_25; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_26; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_27; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_28; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_29; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_30; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_31; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_32; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_33; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_34; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_35; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_36; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_37; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_38; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_39; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_40; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_41; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_42; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_43; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_44; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_45; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_46; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_47; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_48; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_49; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_50; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_51; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_52; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_53; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_54; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_55; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_56; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_57; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_58; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_59; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_60; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_61; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_62; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_63; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_64; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_65; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_66; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_67; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_68; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_69; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_70; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_71; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_72; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_73; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_74; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_75; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_76; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_77; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_78; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_79; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_80; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_81; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_82; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_83; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_84; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_85; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_86; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_87; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_88; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_89; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_90; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_91; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_92; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_93; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_94; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_95; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_96; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_97; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_98; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_99; // @[PEArray.scala 40:21]
  reg [2:0] state; // @[PEArray.scala 100:22]
  wire  _T_3 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_12 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_16 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_22 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_31 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_41 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_342 = _T_41 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 231:12 PEArray.scala 32:8]
  wire  _GEN_349 = _T_31 ? 1'h0 : _GEN_342; // @[Conditional.scala 39:67 PEArray.scala 208:12]
  wire  _GEN_459 = _T_22 | _GEN_349; // @[Conditional.scala 39:67 PEArray.scala 32:8]
  wire  _GEN_463 = _T_16 ? 1'h0 : _GEN_459; // @[Conditional.scala 39:67]
  wire  _GEN_572 = _T_12 | _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 149:12]
  wire  sel1 = _T_3 | _GEN_572; // @[Conditional.scala 40:58 PEArray.scala 108:12]
  wire [15:0] MAC_out = FP16MAC_io_out; // @[PEArray.scala 47:21 PEArray.scala 85:11]
  wire  _GEN_465 = _T_16 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 177:12]
  wire  _GEN_580 = _T_12 | _GEN_465; // @[Conditional.scala 39:67 PEArray.scala 34:8]
  wire  sel3 = _T_3 | _GEN_580; // @[Conditional.scala 40:58 PEArray.scala 110:12]
  wire [1:0] _GEN_344 = _T_41 ? 2'h2 : 2'h0; // @[Conditional.scala 39:67 PEArray.scala 233:12 PEArray.scala 35:8]
  wire [1:0] _GEN_351 = _T_31 ? 2'h2 : _GEN_344; // @[Conditional.scala 39:67 PEArray.scala 210:12]
  wire [1:0] _GEN_461 = _T_22 ? 2'h0 : _GEN_351; // @[Conditional.scala 39:67 PEArray.scala 35:8]
  wire [1:0] _GEN_466 = _T_16 ? 2'h0 : _GEN_461; // @[Conditional.scala 39:67 PEArray.scala 178:12]
  wire [1:0] _GEN_574 = _T_12 ? 2'h1 : _GEN_466; // @[Conditional.scala 39:67]
  wire [1:0] sel4 = _T_3 ? 2'h0 : _GEN_574; // @[Conditional.scala 40:58 PEArray.scala 111:12]
  wire [15:0] _GEN_3 = sel4 == 2'h2 ? io_FromL1 : 16'h0; // @[PEArray.scala 65:28 PEArray.scala 66:15 PEArray.scala 69:15]
  wire [15:0] _GEN_4 = sel4 == 2'h1 ? io_FromAbovePE : _GEN_3; // @[PEArray.scala 62:28 PEArray.scala 63:15]
  wire [15:0] mux4out = sel4 == 2'h0 ? 16'h0 : _GEN_4; // @[PEArray.scala 59:22 PEArray.scala 60:13]
  wire [15:0] _GEN_7 = 6'h1 == L0Index ? L0Memory_1 : L0Memory_0; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_8 = 6'h2 == L0Index ? L0Memory_2 : _GEN_7; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_9 = 6'h3 == L0Index ? L0Memory_3 : _GEN_8; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_10 = 6'h4 == L0Index ? L0Memory_4 : _GEN_9; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_11 = 6'h5 == L0Index ? L0Memory_5 : _GEN_10; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_12 = 6'h6 == L0Index ? L0Memory_6 : _GEN_11; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_13 = 6'h7 == L0Index ? L0Memory_7 : _GEN_12; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_14 = 6'h8 == L0Index ? L0Memory_8 : _GEN_13; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_15 = 6'h9 == L0Index ? L0Memory_9 : _GEN_14; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_16 = 6'ha == L0Index ? L0Memory_10 : _GEN_15; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_17 = 6'hb == L0Index ? L0Memory_11 : _GEN_16; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_18 = 6'hc == L0Index ? L0Memory_12 : _GEN_17; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_19 = 6'hd == L0Index ? L0Memory_13 : _GEN_18; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_20 = 6'he == L0Index ? L0Memory_14 : _GEN_19; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_21 = 6'hf == L0Index ? L0Memory_15 : _GEN_20; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_22 = 6'h10 == L0Index ? L0Memory_16 : _GEN_21; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_23 = 6'h11 == L0Index ? L0Memory_17 : _GEN_22; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_24 = 6'h12 == L0Index ? L0Memory_18 : _GEN_23; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_25 = 6'h13 == L0Index ? L0Memory_19 : _GEN_24; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_26 = 6'h14 == L0Index ? L0Memory_20 : _GEN_25; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_27 = 6'h15 == L0Index ? L0Memory_21 : _GEN_26; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_28 = 6'h16 == L0Index ? L0Memory_22 : _GEN_27; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_29 = 6'h17 == L0Index ? L0Memory_23 : _GEN_28; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_30 = 6'h18 == L0Index ? L0Memory_24 : _GEN_29; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_31 = 6'h19 == L0Index ? L0Memory_25 : _GEN_30; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_32 = 6'h1a == L0Index ? L0Memory_26 : _GEN_31; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_33 = 6'h1b == L0Index ? L0Memory_27 : _GEN_32; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_34 = 6'h1c == L0Index ? L0Memory_28 : _GEN_33; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_35 = 6'h1d == L0Index ? L0Memory_29 : _GEN_34; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_36 = 6'h1e == L0Index ? L0Memory_30 : _GEN_35; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_37 = 6'h1f == L0Index ? L0Memory_31 : _GEN_36; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_38 = 6'h20 == L0Index ? L0Memory_32 : _GEN_37; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_39 = 6'h21 == L0Index ? L0Memory_33 : _GEN_38; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_40 = 6'h22 == L0Index ? L0Memory_34 : _GEN_39; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_41 = 6'h23 == L0Index ? L0Memory_35 : _GEN_40; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_42 = 6'h24 == L0Index ? L0Memory_36 : _GEN_41; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_43 = 6'h25 == L0Index ? L0Memory_37 : _GEN_42; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_44 = 6'h26 == L0Index ? L0Memory_38 : _GEN_43; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_45 = 6'h27 == L0Index ? L0Memory_39 : _GEN_44; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_46 = 6'h28 == L0Index ? L0Memory_40 : _GEN_45; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_47 = 6'h29 == L0Index ? L0Memory_41 : _GEN_46; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_48 = 6'h2a == L0Index ? L0Memory_42 : _GEN_47; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_49 = 6'h2b == L0Index ? L0Memory_43 : _GEN_48; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_50 = 6'h2c == L0Index ? L0Memory_44 : _GEN_49; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_51 = 6'h2d == L0Index ? L0Memory_45 : _GEN_50; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_52 = 6'h2e == L0Index ? L0Memory_46 : _GEN_51; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_53 = 6'h2f == L0Index ? L0Memory_47 : _GEN_52; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_54 = 6'h30 == L0Index ? L0Memory_48 : _GEN_53; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_55 = 6'h31 == L0Index ? L0Memory_49 : _GEN_54; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_56 = 6'h32 == L0Index ? L0Memory_50 : _GEN_55; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_57 = 6'h33 == L0Index ? L0Memory_51 : _GEN_56; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_58 = 6'h34 == L0Index ? L0Memory_52 : _GEN_57; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_59 = 6'h35 == L0Index ? L0Memory_53 : _GEN_58; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_60 = 6'h36 == L0Index ? L0Memory_54 : _GEN_59; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_61 = 6'h37 == L0Index ? L0Memory_55 : _GEN_60; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_62 = 6'h38 == L0Index ? L0Memory_56 : _GEN_61; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_63 = 6'h39 == L0Index ? L0Memory_57 : _GEN_62; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_64 = 6'h3a == L0Index ? L0Memory_58 : _GEN_63; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_65 = 6'h3b == L0Index ? L0Memory_59 : _GEN_64; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_66 = 6'h3c == L0Index ? L0Memory_60 : _GEN_65; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_67 = 6'h3d == L0Index ? L0Memory_61 : _GEN_66; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_68 = 6'h3e == L0Index ? L0Memory_62 : _GEN_67; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_69 = 6'h3f == L0Index ? L0Memory_63 : _GEN_68; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [6:0] _GEN_793 = {{1'd0}, L0Index}; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_70 = 7'h40 == _GEN_793 ? L0Memory_64 : _GEN_69; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_71 = 7'h41 == _GEN_793 ? L0Memory_65 : _GEN_70; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_72 = 7'h42 == _GEN_793 ? L0Memory_66 : _GEN_71; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_73 = 7'h43 == _GEN_793 ? L0Memory_67 : _GEN_72; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_74 = 7'h44 == _GEN_793 ? L0Memory_68 : _GEN_73; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_75 = 7'h45 == _GEN_793 ? L0Memory_69 : _GEN_74; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_76 = 7'h46 == _GEN_793 ? L0Memory_70 : _GEN_75; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_77 = 7'h47 == _GEN_793 ? L0Memory_71 : _GEN_76; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_78 = 7'h48 == _GEN_793 ? L0Memory_72 : _GEN_77; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_79 = 7'h49 == _GEN_793 ? L0Memory_73 : _GEN_78; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_80 = 7'h4a == _GEN_793 ? L0Memory_74 : _GEN_79; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_81 = 7'h4b == _GEN_793 ? L0Memory_75 : _GEN_80; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_82 = 7'h4c == _GEN_793 ? L0Memory_76 : _GEN_81; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_83 = 7'h4d == _GEN_793 ? L0Memory_77 : _GEN_82; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_84 = 7'h4e == _GEN_793 ? L0Memory_78 : _GEN_83; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_85 = 7'h4f == _GEN_793 ? L0Memory_79 : _GEN_84; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_86 = 7'h50 == _GEN_793 ? L0Memory_80 : _GEN_85; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_87 = 7'h51 == _GEN_793 ? L0Memory_81 : _GEN_86; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_88 = 7'h52 == _GEN_793 ? L0Memory_82 : _GEN_87; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_89 = 7'h53 == _GEN_793 ? L0Memory_83 : _GEN_88; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_90 = 7'h54 == _GEN_793 ? L0Memory_84 : _GEN_89; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_91 = 7'h55 == _GEN_793 ? L0Memory_85 : _GEN_90; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_92 = 7'h56 == _GEN_793 ? L0Memory_86 : _GEN_91; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_93 = 7'h57 == _GEN_793 ? L0Memory_87 : _GEN_92; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_94 = 7'h58 == _GEN_793 ? L0Memory_88 : _GEN_93; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_95 = 7'h59 == _GEN_793 ? L0Memory_89 : _GEN_94; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_96 = 7'h5a == _GEN_793 ? L0Memory_90 : _GEN_95; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_97 = 7'h5b == _GEN_793 ? L0Memory_91 : _GEN_96; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_98 = 7'h5c == _GEN_793 ? L0Memory_92 : _GEN_97; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_99 = 7'h5d == _GEN_793 ? L0Memory_93 : _GEN_98; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_100 = 7'h5e == _GEN_793 ? L0Memory_94 : _GEN_99; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_101 = 7'h5f == _GEN_793 ? L0Memory_95 : _GEN_100; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_102 = 7'h60 == _GEN_793 ? L0Memory_96 : _GEN_101; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_103 = 7'h61 == _GEN_793 ? L0Memory_97 : _GEN_102; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_104 = 7'h62 == _GEN_793 ? L0Memory_98 : _GEN_103; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_105 = 7'h63 == _GEN_793 ? L0Memory_99 : _GEN_104; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire  _GEN_575 = _T_12 ? 1'h0 : _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 157:12]
  wire  sel5 = _T_3 ? 1'h0 : _GEN_575; // @[Conditional.scala 40:58 PEArray.scala 112:12]
  reg [15:0] mux2out_reg; // @[PEArray.scala 90:28]
  reg [15:0] mux3out_reg; // @[PEArray.scala 91:28]
  reg [9:0] count; // @[PEArray.scala 101:22]
  reg [5:0] GRU_out_width; // @[PEArray.scala 104:26]
  wire [7:0] _GEN_118 = io_control_signal_mask[9] ? 8'h0 : {{2'd0}, GRU_out_width}; // @[PEArray.scala 116:57 PEArray.scala 145:23 PEArray.scala 104:26]
  wire [9:0] _count_T_1 = count + 10'h1; // @[PEArray.scala 162:24]
  wire [9:0] _GEN_120 = count != 10'h33 ? _count_T_1 : count; // @[PEArray.scala 161:27 PEArray.scala 162:15 PEArray.scala 101:22]
  wire [9:0] _GEN_124 = count != 10'h188 ? _count_T_1 : count; // @[PEArray.scala 183:28 PEArray.scala 184:15 PEArray.scala 101:22]
  wire [9:0] _GEN_125 = count == 10'h188 ? 10'h0 : _GEN_124; // @[PEArray.scala 186:28 PEArray.scala 187:15]
  wire [2:0] _GEN_126 = count == 10'h188 ? 3'h0 : state; // @[PEArray.scala 186:28 PEArray.scala 188:15 PEArray.scala 100:22]
  wire [9:0] _GEN_127 = count != 10'h0 ? _count_T_1 : count; // @[PEArray.scala 192:32 PEArray.scala 193:15 PEArray.scala 101:22]
  wire  _T_24 = count == 10'h0; // @[PEArray.scala 195:18]
  wire [5:0] _GEN_128 = count == 10'h0 ? 6'h0 : L0Index; // @[PEArray.scala 195:26 PEArray.scala 196:17 PEArray.scala 39:24]
  wire [9:0] _T_27 = 10'h0 - 10'h1; // @[PEArray.scala 198:51]
  wire [15:0] _GEN_129 = 6'h0 == L0Index ? io_FromL1 : L0Memory_0; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_130 = 6'h1 == L0Index ? io_FromL1 : L0Memory_1; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_131 = 6'h2 == L0Index ? io_FromL1 : L0Memory_2; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_132 = 6'h3 == L0Index ? io_FromL1 : L0Memory_3; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_133 = 6'h4 == L0Index ? io_FromL1 : L0Memory_4; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_134 = 6'h5 == L0Index ? io_FromL1 : L0Memory_5; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_135 = 6'h6 == L0Index ? io_FromL1 : L0Memory_6; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_136 = 6'h7 == L0Index ? io_FromL1 : L0Memory_7; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_137 = 6'h8 == L0Index ? io_FromL1 : L0Memory_8; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_138 = 6'h9 == L0Index ? io_FromL1 : L0Memory_9; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_139 = 6'ha == L0Index ? io_FromL1 : L0Memory_10; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_140 = 6'hb == L0Index ? io_FromL1 : L0Memory_11; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_141 = 6'hc == L0Index ? io_FromL1 : L0Memory_12; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_142 = 6'hd == L0Index ? io_FromL1 : L0Memory_13; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_143 = 6'he == L0Index ? io_FromL1 : L0Memory_14; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_144 = 6'hf == L0Index ? io_FromL1 : L0Memory_15; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_145 = 6'h10 == L0Index ? io_FromL1 : L0Memory_16; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_146 = 6'h11 == L0Index ? io_FromL1 : L0Memory_17; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_147 = 6'h12 == L0Index ? io_FromL1 : L0Memory_18; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_148 = 6'h13 == L0Index ? io_FromL1 : L0Memory_19; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_149 = 6'h14 == L0Index ? io_FromL1 : L0Memory_20; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_150 = 6'h15 == L0Index ? io_FromL1 : L0Memory_21; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_151 = 6'h16 == L0Index ? io_FromL1 : L0Memory_22; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_152 = 6'h17 == L0Index ? io_FromL1 : L0Memory_23; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_153 = 6'h18 == L0Index ? io_FromL1 : L0Memory_24; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_154 = 6'h19 == L0Index ? io_FromL1 : L0Memory_25; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_155 = 6'h1a == L0Index ? io_FromL1 : L0Memory_26; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_156 = 6'h1b == L0Index ? io_FromL1 : L0Memory_27; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_157 = 6'h1c == L0Index ? io_FromL1 : L0Memory_28; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_158 = 6'h1d == L0Index ? io_FromL1 : L0Memory_29; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_159 = 6'h1e == L0Index ? io_FromL1 : L0Memory_30; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_160 = 6'h1f == L0Index ? io_FromL1 : L0Memory_31; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_161 = 6'h20 == L0Index ? io_FromL1 : L0Memory_32; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_162 = 6'h21 == L0Index ? io_FromL1 : L0Memory_33; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_163 = 6'h22 == L0Index ? io_FromL1 : L0Memory_34; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_164 = 6'h23 == L0Index ? io_FromL1 : L0Memory_35; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_165 = 6'h24 == L0Index ? io_FromL1 : L0Memory_36; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_166 = 6'h25 == L0Index ? io_FromL1 : L0Memory_37; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_167 = 6'h26 == L0Index ? io_FromL1 : L0Memory_38; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_168 = 6'h27 == L0Index ? io_FromL1 : L0Memory_39; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_169 = 6'h28 == L0Index ? io_FromL1 : L0Memory_40; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_170 = 6'h29 == L0Index ? io_FromL1 : L0Memory_41; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_171 = 6'h2a == L0Index ? io_FromL1 : L0Memory_42; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_172 = 6'h2b == L0Index ? io_FromL1 : L0Memory_43; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_173 = 6'h2c == L0Index ? io_FromL1 : L0Memory_44; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_174 = 6'h2d == L0Index ? io_FromL1 : L0Memory_45; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_175 = 6'h2e == L0Index ? io_FromL1 : L0Memory_46; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_176 = 6'h2f == L0Index ? io_FromL1 : L0Memory_47; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_177 = 6'h30 == L0Index ? io_FromL1 : L0Memory_48; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_178 = 6'h31 == L0Index ? io_FromL1 : L0Memory_49; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_179 = 6'h32 == L0Index ? io_FromL1 : L0Memory_50; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_180 = 6'h33 == L0Index ? io_FromL1 : L0Memory_51; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_181 = 6'h34 == L0Index ? io_FromL1 : L0Memory_52; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_182 = 6'h35 == L0Index ? io_FromL1 : L0Memory_53; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_183 = 6'h36 == L0Index ? io_FromL1 : L0Memory_54; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_184 = 6'h37 == L0Index ? io_FromL1 : L0Memory_55; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_185 = 6'h38 == L0Index ? io_FromL1 : L0Memory_56; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_186 = 6'h39 == L0Index ? io_FromL1 : L0Memory_57; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_187 = 6'h3a == L0Index ? io_FromL1 : L0Memory_58; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_188 = 6'h3b == L0Index ? io_FromL1 : L0Memory_59; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_189 = 6'h3c == L0Index ? io_FromL1 : L0Memory_60; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_190 = 6'h3d == L0Index ? io_FromL1 : L0Memory_61; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_191 = 6'h3e == L0Index ? io_FromL1 : L0Memory_62; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_192 = 6'h3f == L0Index ? io_FromL1 : L0Memory_63; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_193 = 7'h40 == _GEN_793 ? io_FromL1 : L0Memory_64; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_194 = 7'h41 == _GEN_793 ? io_FromL1 : L0Memory_65; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_195 = 7'h42 == _GEN_793 ? io_FromL1 : L0Memory_66; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_196 = 7'h43 == _GEN_793 ? io_FromL1 : L0Memory_67; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_197 = 7'h44 == _GEN_793 ? io_FromL1 : L0Memory_68; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_198 = 7'h45 == _GEN_793 ? io_FromL1 : L0Memory_69; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_199 = 7'h46 == _GEN_793 ? io_FromL1 : L0Memory_70; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_200 = 7'h47 == _GEN_793 ? io_FromL1 : L0Memory_71; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_201 = 7'h48 == _GEN_793 ? io_FromL1 : L0Memory_72; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_202 = 7'h49 == _GEN_793 ? io_FromL1 : L0Memory_73; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_203 = 7'h4a == _GEN_793 ? io_FromL1 : L0Memory_74; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_204 = 7'h4b == _GEN_793 ? io_FromL1 : L0Memory_75; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_205 = 7'h4c == _GEN_793 ? io_FromL1 : L0Memory_76; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_206 = 7'h4d == _GEN_793 ? io_FromL1 : L0Memory_77; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_207 = 7'h4e == _GEN_793 ? io_FromL1 : L0Memory_78; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_208 = 7'h4f == _GEN_793 ? io_FromL1 : L0Memory_79; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_209 = 7'h50 == _GEN_793 ? io_FromL1 : L0Memory_80; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_210 = 7'h51 == _GEN_793 ? io_FromL1 : L0Memory_81; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_211 = 7'h52 == _GEN_793 ? io_FromL1 : L0Memory_82; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_212 = 7'h53 == _GEN_793 ? io_FromL1 : L0Memory_83; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_213 = 7'h54 == _GEN_793 ? io_FromL1 : L0Memory_84; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_214 = 7'h55 == _GEN_793 ? io_FromL1 : L0Memory_85; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_215 = 7'h56 == _GEN_793 ? io_FromL1 : L0Memory_86; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_216 = 7'h57 == _GEN_793 ? io_FromL1 : L0Memory_87; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_217 = 7'h58 == _GEN_793 ? io_FromL1 : L0Memory_88; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_218 = 7'h59 == _GEN_793 ? io_FromL1 : L0Memory_89; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_219 = 7'h5a == _GEN_793 ? io_FromL1 : L0Memory_90; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_220 = 7'h5b == _GEN_793 ? io_FromL1 : L0Memory_91; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_221 = 7'h5c == _GEN_793 ? io_FromL1 : L0Memory_92; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_222 = 7'h5d == _GEN_793 ? io_FromL1 : L0Memory_93; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_223 = 7'h5e == _GEN_793 ? io_FromL1 : L0Memory_94; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_224 = 7'h5f == _GEN_793 ? io_FromL1 : L0Memory_95; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_225 = 7'h60 == _GEN_793 ? io_FromL1 : L0Memory_96; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_226 = 7'h61 == _GEN_793 ? io_FromL1 : L0Memory_97; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_227 = 7'h62 == _GEN_793 ? io_FromL1 : L0Memory_98; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_228 = 7'h63 == _GEN_793 ? io_FromL1 : L0Memory_99; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [5:0] _L0Index_T_2 = L0Index + 6'h1; // @[PEArray.scala 200:28]
  wire [15:0] _GEN_229 = count >= 10'h1 & count <= _T_27 ? _GEN_129 : L0Memory_0; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_230 = count >= 10'h1 & count <= _T_27 ? _GEN_130 : L0Memory_1; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_231 = count >= 10'h1 & count <= _T_27 ? _GEN_131 : L0Memory_2; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_232 = count >= 10'h1 & count <= _T_27 ? _GEN_132 : L0Memory_3; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_233 = count >= 10'h1 & count <= _T_27 ? _GEN_133 : L0Memory_4; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_234 = count >= 10'h1 & count <= _T_27 ? _GEN_134 : L0Memory_5; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_235 = count >= 10'h1 & count <= _T_27 ? _GEN_135 : L0Memory_6; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_236 = count >= 10'h1 & count <= _T_27 ? _GEN_136 : L0Memory_7; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_237 = count >= 10'h1 & count <= _T_27 ? _GEN_137 : L0Memory_8; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_238 = count >= 10'h1 & count <= _T_27 ? _GEN_138 : L0Memory_9; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_239 = count >= 10'h1 & count <= _T_27 ? _GEN_139 : L0Memory_10; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_240 = count >= 10'h1 & count <= _T_27 ? _GEN_140 : L0Memory_11; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_241 = count >= 10'h1 & count <= _T_27 ? _GEN_141 : L0Memory_12; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_242 = count >= 10'h1 & count <= _T_27 ? _GEN_142 : L0Memory_13; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_243 = count >= 10'h1 & count <= _T_27 ? _GEN_143 : L0Memory_14; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_244 = count >= 10'h1 & count <= _T_27 ? _GEN_144 : L0Memory_15; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_245 = count >= 10'h1 & count <= _T_27 ? _GEN_145 : L0Memory_16; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_246 = count >= 10'h1 & count <= _T_27 ? _GEN_146 : L0Memory_17; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_247 = count >= 10'h1 & count <= _T_27 ? _GEN_147 : L0Memory_18; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_248 = count >= 10'h1 & count <= _T_27 ? _GEN_148 : L0Memory_19; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_249 = count >= 10'h1 & count <= _T_27 ? _GEN_149 : L0Memory_20; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_250 = count >= 10'h1 & count <= _T_27 ? _GEN_150 : L0Memory_21; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_251 = count >= 10'h1 & count <= _T_27 ? _GEN_151 : L0Memory_22; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_252 = count >= 10'h1 & count <= _T_27 ? _GEN_152 : L0Memory_23; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_253 = count >= 10'h1 & count <= _T_27 ? _GEN_153 : L0Memory_24; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_254 = count >= 10'h1 & count <= _T_27 ? _GEN_154 : L0Memory_25; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_255 = count >= 10'h1 & count <= _T_27 ? _GEN_155 : L0Memory_26; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_256 = count >= 10'h1 & count <= _T_27 ? _GEN_156 : L0Memory_27; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_257 = count >= 10'h1 & count <= _T_27 ? _GEN_157 : L0Memory_28; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_258 = count >= 10'h1 & count <= _T_27 ? _GEN_158 : L0Memory_29; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_259 = count >= 10'h1 & count <= _T_27 ? _GEN_159 : L0Memory_30; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_260 = count >= 10'h1 & count <= _T_27 ? _GEN_160 : L0Memory_31; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_261 = count >= 10'h1 & count <= _T_27 ? _GEN_161 : L0Memory_32; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_262 = count >= 10'h1 & count <= _T_27 ? _GEN_162 : L0Memory_33; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_263 = count >= 10'h1 & count <= _T_27 ? _GEN_163 : L0Memory_34; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_264 = count >= 10'h1 & count <= _T_27 ? _GEN_164 : L0Memory_35; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_265 = count >= 10'h1 & count <= _T_27 ? _GEN_165 : L0Memory_36; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_266 = count >= 10'h1 & count <= _T_27 ? _GEN_166 : L0Memory_37; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_267 = count >= 10'h1 & count <= _T_27 ? _GEN_167 : L0Memory_38; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_268 = count >= 10'h1 & count <= _T_27 ? _GEN_168 : L0Memory_39; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_269 = count >= 10'h1 & count <= _T_27 ? _GEN_169 : L0Memory_40; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_270 = count >= 10'h1 & count <= _T_27 ? _GEN_170 : L0Memory_41; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_271 = count >= 10'h1 & count <= _T_27 ? _GEN_171 : L0Memory_42; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_272 = count >= 10'h1 & count <= _T_27 ? _GEN_172 : L0Memory_43; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_273 = count >= 10'h1 & count <= _T_27 ? _GEN_173 : L0Memory_44; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_274 = count >= 10'h1 & count <= _T_27 ? _GEN_174 : L0Memory_45; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_275 = count >= 10'h1 & count <= _T_27 ? _GEN_175 : L0Memory_46; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_276 = count >= 10'h1 & count <= _T_27 ? _GEN_176 : L0Memory_47; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_277 = count >= 10'h1 & count <= _T_27 ? _GEN_177 : L0Memory_48; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_278 = count >= 10'h1 & count <= _T_27 ? _GEN_178 : L0Memory_49; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_279 = count >= 10'h1 & count <= _T_27 ? _GEN_179 : L0Memory_50; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_280 = count >= 10'h1 & count <= _T_27 ? _GEN_180 : L0Memory_51; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_281 = count >= 10'h1 & count <= _T_27 ? _GEN_181 : L0Memory_52; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_282 = count >= 10'h1 & count <= _T_27 ? _GEN_182 : L0Memory_53; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_283 = count >= 10'h1 & count <= _T_27 ? _GEN_183 : L0Memory_54; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_284 = count >= 10'h1 & count <= _T_27 ? _GEN_184 : L0Memory_55; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_285 = count >= 10'h1 & count <= _T_27 ? _GEN_185 : L0Memory_56; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_286 = count >= 10'h1 & count <= _T_27 ? _GEN_186 : L0Memory_57; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_287 = count >= 10'h1 & count <= _T_27 ? _GEN_187 : L0Memory_58; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_288 = count >= 10'h1 & count <= _T_27 ? _GEN_188 : L0Memory_59; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_289 = count >= 10'h1 & count <= _T_27 ? _GEN_189 : L0Memory_60; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_290 = count >= 10'h1 & count <= _T_27 ? _GEN_190 : L0Memory_61; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_291 = count >= 10'h1 & count <= _T_27 ? _GEN_191 : L0Memory_62; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_292 = count >= 10'h1 & count <= _T_27 ? _GEN_192 : L0Memory_63; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_293 = count >= 10'h1 & count <= _T_27 ? _GEN_193 : L0Memory_64; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_294 = count >= 10'h1 & count <= _T_27 ? _GEN_194 : L0Memory_65; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_295 = count >= 10'h1 & count <= _T_27 ? _GEN_195 : L0Memory_66; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_296 = count >= 10'h1 & count <= _T_27 ? _GEN_196 : L0Memory_67; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_297 = count >= 10'h1 & count <= _T_27 ? _GEN_197 : L0Memory_68; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_298 = count >= 10'h1 & count <= _T_27 ? _GEN_198 : L0Memory_69; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_299 = count >= 10'h1 & count <= _T_27 ? _GEN_199 : L0Memory_70; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_300 = count >= 10'h1 & count <= _T_27 ? _GEN_200 : L0Memory_71; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_301 = count >= 10'h1 & count <= _T_27 ? _GEN_201 : L0Memory_72; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_302 = count >= 10'h1 & count <= _T_27 ? _GEN_202 : L0Memory_73; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_303 = count >= 10'h1 & count <= _T_27 ? _GEN_203 : L0Memory_74; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_304 = count >= 10'h1 & count <= _T_27 ? _GEN_204 : L0Memory_75; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_305 = count >= 10'h1 & count <= _T_27 ? _GEN_205 : L0Memory_76; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_306 = count >= 10'h1 & count <= _T_27 ? _GEN_206 : L0Memory_77; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_307 = count >= 10'h1 & count <= _T_27 ? _GEN_207 : L0Memory_78; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_308 = count >= 10'h1 & count <= _T_27 ? _GEN_208 : L0Memory_79; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_309 = count >= 10'h1 & count <= _T_27 ? _GEN_209 : L0Memory_80; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_310 = count >= 10'h1 & count <= _T_27 ? _GEN_210 : L0Memory_81; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_311 = count >= 10'h1 & count <= _T_27 ? _GEN_211 : L0Memory_82; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_312 = count >= 10'h1 & count <= _T_27 ? _GEN_212 : L0Memory_83; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_313 = count >= 10'h1 & count <= _T_27 ? _GEN_213 : L0Memory_84; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_314 = count >= 10'h1 & count <= _T_27 ? _GEN_214 : L0Memory_85; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_315 = count >= 10'h1 & count <= _T_27 ? _GEN_215 : L0Memory_86; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_316 = count >= 10'h1 & count <= _T_27 ? _GEN_216 : L0Memory_87; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_317 = count >= 10'h1 & count <= _T_27 ? _GEN_217 : L0Memory_88; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_318 = count >= 10'h1 & count <= _T_27 ? _GEN_218 : L0Memory_89; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_319 = count >= 10'h1 & count <= _T_27 ? _GEN_219 : L0Memory_90; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_320 = count >= 10'h1 & count <= _T_27 ? _GEN_220 : L0Memory_91; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_321 = count >= 10'h1 & count <= _T_27 ? _GEN_221 : L0Memory_92; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_322 = count >= 10'h1 & count <= _T_27 ? _GEN_222 : L0Memory_93; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_323 = count >= 10'h1 & count <= _T_27 ? _GEN_223 : L0Memory_94; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_324 = count >= 10'h1 & count <= _T_27 ? _GEN_224 : L0Memory_95; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_325 = count >= 10'h1 & count <= _T_27 ? _GEN_225 : L0Memory_96; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_326 = count >= 10'h1 & count <= _T_27 ? _GEN_226 : L0Memory_97; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_327 = count >= 10'h1 & count <= _T_27 ? _GEN_227 : L0Memory_98; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_328 = count >= 10'h1 & count <= _T_27 ? _GEN_228 : L0Memory_99; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [5:0] _GEN_329 = count >= 10'h1 & count <= _T_27 ? _L0Index_T_2 : _GEN_128; // @[PEArray.scala 198:59 PEArray.scala 200:17]
  wire [9:0] _GEN_330 = _T_24 ? 10'h0 : _GEN_127; // @[PEArray.scala 202:32 PEArray.scala 203:15]
  wire [2:0] _GEN_331 = _T_24 ? 3'h0 : state; // @[PEArray.scala 202:32 PEArray.scala 204:15 PEArray.scala 100:22]
  wire [9:0] _GEN_865 = {{4'd0}, GRU_out_width}; // @[PEArray.scala 220:19]
  wire [9:0] _GEN_0 = count % _GEN_865; // @[PEArray.scala 220:19]
  wire [5:0] _T_36 = _GEN_0[5:0]; // @[PEArray.scala 220:19]
  wire [5:0] _T_38 = GRU_out_width - 6'h1; // @[PEArray.scala 220:55]
  wire [5:0] _GEN_334 = _T_36 == _T_38 ? _L0Index_T_2 : 6'h0; // @[PEArray.scala 220:62 PEArray.scala 221:17 PEArray.scala 214:15]
  wire [5:0] _GEN_346 = _T_41 ? _GEN_334 : L0Index; // @[Conditional.scala 39:67 PEArray.scala 39:24]
  wire [9:0] _GEN_347 = _T_41 ? _GEN_330 : count; // @[Conditional.scala 39:67 PEArray.scala 101:22]
  wire [2:0] _GEN_348 = _T_41 ? _GEN_331 : state; // @[Conditional.scala 39:67 PEArray.scala 100:22]
  wire [5:0] _GEN_353 = _T_31 ? _GEN_334 : _GEN_346; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_354 = _T_31 ? _GEN_330 : _GEN_347; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_355 = _T_31 ? _GEN_331 : _GEN_348; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_356 = _T_22 ? _GEN_330 : _GEN_354; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_357 = _T_22 ? _GEN_329 : _GEN_353; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_458 = _T_22 ? _GEN_331 : _GEN_355; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_690 = _T_3 ? _GEN_118 : {{2'd0}, GRU_out_width}; // @[Conditional.scala 40:58 PEArray.scala 104:26]
  FP16MulAdder FP16MAC ( // @[PEArray.scala 72:23]
    .io_a(FP16MAC_io_a),
    .io_b(FP16MAC_io_b),
    .io_c(FP16MAC_io_c),
    .io_out(FP16MAC_io_out)
  );
  assign io_ToRightPE = mux3out_reg; // @[PEArray.scala 95:16]
  assign io_ToBelowPE = mux2out_reg; // @[PEArray.scala 94:16]
  assign FP16MAC_io_a = sel1 ? io_FromL1 : io_FromLeftPE; // @[PEArray.scala 50:14 PEArray.scala 50:23 PEArray.scala 51:24]
  assign FP16MAC_io_b = sel5 ? mux4out : _GEN_105; // @[PEArray.scala 77:13 PEArray.scala 78:18 PEArray.scala 81:18]
  assign FP16MAC_io_c = sel5 ? _GEN_105 : mux4out; // @[PEArray.scala 77:13 PEArray.scala 79:18 PEArray.scala 82:18]
  always @(posedge clock) begin
    if (reset) begin // @[PEArray.scala 39:24]
      L0Index <= 6'h0; // @[PEArray.scala 39:24]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h1; // @[PEArray.scala 159:15]
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h5; // @[PEArray.scala 181:15]
      end else begin
        L0Index <= _GEN_357;
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_0 <= _GEN_229;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_1 <= _GEN_230;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_2 <= _GEN_231;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_3 <= _GEN_232;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_4 <= _GEN_233;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_5 <= _GEN_234;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_6 <= _GEN_235;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_7 <= _GEN_236;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_8 <= _GEN_237;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_9 <= _GEN_238;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_10 <= _GEN_239;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_11 <= _GEN_240;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_12 <= _GEN_241;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_13 <= _GEN_242;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_14 <= _GEN_243;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_15 <= _GEN_244;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_16 <= _GEN_245;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_17 <= _GEN_246;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_18 <= _GEN_247;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_19 <= _GEN_248;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_20 <= _GEN_249;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_21 <= _GEN_250;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_22 <= _GEN_251;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_23 <= _GEN_252;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_24 <= _GEN_253;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_25 <= _GEN_254;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_26 <= _GEN_255;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_27 <= _GEN_256;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_28 <= _GEN_257;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_29 <= _GEN_258;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_30 <= _GEN_259;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_31 <= _GEN_260;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_32 <= _GEN_261;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_33 <= _GEN_262;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_34 <= _GEN_263;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_35 <= _GEN_264;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_36 <= _GEN_265;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_37 <= _GEN_266;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_38 <= _GEN_267;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_39 <= _GEN_268;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_40 <= _GEN_269;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_41 <= _GEN_270;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_42 <= _GEN_271;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_43 <= _GEN_272;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_44 <= _GEN_273;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_45 <= _GEN_274;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_46 <= _GEN_275;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_47 <= _GEN_276;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_48 <= _GEN_277;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_49 <= _GEN_278;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_50 <= _GEN_279;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_51 <= _GEN_280;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_52 <= _GEN_281;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_53 <= _GEN_282;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_54 <= _GEN_283;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_55 <= _GEN_284;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_56 <= _GEN_285;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_57 <= _GEN_286;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_58 <= _GEN_287;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_59 <= _GEN_288;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_60 <= _GEN_289;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_61 <= _GEN_290;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_62 <= _GEN_291;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_63 <= _GEN_292;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_64 <= _GEN_293;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_65 <= _GEN_294;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_66 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_67 <= _GEN_296;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_68 <= _GEN_297;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_69 <= _GEN_298;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_70 <= _GEN_299;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_71 <= _GEN_300;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_72 <= _GEN_301;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_73 <= _GEN_302;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_74 <= _GEN_303;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_75 <= _GEN_304;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_76 <= _GEN_305;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_77 <= _GEN_306;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_78 <= _GEN_307;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_79 <= _GEN_308;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_80 <= _GEN_309;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_81 <= _GEN_310;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_82 <= _GEN_311;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_83 <= _GEN_312;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_84 <= _GEN_313;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_85 <= _GEN_314;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_86 <= _GEN_315;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_87 <= _GEN_316;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_88 <= _GEN_317;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_89 <= _GEN_318;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_90 <= _GEN_319;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_91 <= _GEN_320;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_92 <= _GEN_321;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_93 <= _GEN_322;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_94 <= _GEN_323;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_95 <= _GEN_324;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_96 <= _GEN_325;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_97 <= _GEN_326;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_98 <= _GEN_327;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_99 <= _GEN_328;
          end
        end
      end
    end
    if (reset) begin // @[PEArray.scala 100:22]
      state <= 3'h0; // @[PEArray.scala 100:22]
    end else if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[9]) begin // @[PEArray.scala 116:57]
        state <= 3'h1;
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      if (count == 10'h33) begin // @[PEArray.scala 164:27]
        state <= 3'h0; // @[PEArray.scala 166:15]
      end
    end else if (_T_16) begin // @[Conditional.scala 39:67]
      state <= _GEN_126;
    end else begin
      state <= _GEN_458;
    end
    if (reset) begin // @[PEArray.scala 90:28]
      mux2out_reg <= 16'h0; // @[PEArray.scala 90:28]
    end else begin
      mux2out_reg <= MAC_out; // @[PEArray.scala 90:28]
    end
    if (reset) begin // @[PEArray.scala 91:28]
      mux3out_reg <= 16'h0; // @[PEArray.scala 91:28]
    end else if (sel3) begin // @[PEArray.scala 56:14]
      mux3out_reg <= MAC_out; // @[PEArray.scala 56:23]
    end else if (sel1) begin // @[PEArray.scala 50:14]
      mux3out_reg <= io_FromL1; // @[PEArray.scala 50:23]
    end else begin
      mux3out_reg <= io_FromLeftPE; // @[PEArray.scala 51:24]
    end
    if (reset) begin // @[PEArray.scala 101:22]
      count <= 10'h0; // @[PEArray.scala 101:22]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        if (count == 10'h33) begin // @[PEArray.scala 164:27]
          count <= 10'h0; // @[PEArray.scala 165:15]
        end else begin
          count <= _GEN_120;
        end
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        count <= _GEN_125;
      end else begin
        count <= _GEN_356;
      end
    end
    GRU_out_width <= _GEN_690[5:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  L0Index = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  L0Memory_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  L0Memory_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  L0Memory_2 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  L0Memory_3 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  L0Memory_4 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  L0Memory_5 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  L0Memory_6 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  L0Memory_7 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  L0Memory_8 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  L0Memory_9 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  L0Memory_10 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  L0Memory_11 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  L0Memory_12 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  L0Memory_13 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  L0Memory_14 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  L0Memory_15 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  L0Memory_16 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  L0Memory_17 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  L0Memory_18 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  L0Memory_19 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  L0Memory_20 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  L0Memory_21 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  L0Memory_22 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  L0Memory_23 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  L0Memory_24 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  L0Memory_25 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  L0Memory_26 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  L0Memory_27 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  L0Memory_28 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  L0Memory_29 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  L0Memory_30 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  L0Memory_31 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  L0Memory_32 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  L0Memory_33 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  L0Memory_34 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  L0Memory_35 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  L0Memory_36 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  L0Memory_37 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  L0Memory_38 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  L0Memory_39 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  L0Memory_40 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  L0Memory_41 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  L0Memory_42 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  L0Memory_43 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  L0Memory_44 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  L0Memory_45 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  L0Memory_46 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  L0Memory_47 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  L0Memory_48 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  L0Memory_49 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  L0Memory_50 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  L0Memory_51 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  L0Memory_52 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  L0Memory_53 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  L0Memory_54 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  L0Memory_55 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  L0Memory_56 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  L0Memory_57 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  L0Memory_58 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  L0Memory_59 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  L0Memory_60 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  L0Memory_61 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  L0Memory_62 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  L0Memory_63 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  L0Memory_64 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  L0Memory_65 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  L0Memory_66 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  L0Memory_67 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  L0Memory_68 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  L0Memory_69 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  L0Memory_70 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  L0Memory_71 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  L0Memory_72 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  L0Memory_73 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  L0Memory_74 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  L0Memory_75 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  L0Memory_76 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  L0Memory_77 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  L0Memory_78 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  L0Memory_79 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  L0Memory_80 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  L0Memory_81 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  L0Memory_82 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  L0Memory_83 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  L0Memory_84 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  L0Memory_85 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  L0Memory_86 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  L0Memory_87 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  L0Memory_88 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  L0Memory_89 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  L0Memory_90 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  L0Memory_91 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  L0Memory_92 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  L0Memory_93 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  L0Memory_94 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  L0Memory_95 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  L0Memory_96 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  L0Memory_97 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  L0Memory_98 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  L0Memory_99 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  state = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  mux2out_reg = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  mux3out_reg = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  count = _RAND_104[9:0];
  _RAND_105 = {1{`RANDOM}};
  GRU_out_width = _RAND_105[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PE_8(
  input         clock,
  input         reset,
  input  [15:0] io_FromAbovePE,
  input  [15:0] io_FromLeftPE,
  input  [15:0] io_FromL1,
  input  [2:0]  io_control_signal_control,
  input  [9:0]  io_control_signal_count,
  input  [5:0]  io_control_signal_L0index,
  input  [11:0] io_control_signal_mask,
  input  [7:0]  io_control_signal_gru_out_width,
  output [15:0] io_ToRightPE,
  output [15:0] io_ToBelowPE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] FP16MAC_io_a; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_b; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_c; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_out; // @[PEArray.scala 72:23]
  reg [5:0] L0Index; // @[PEArray.scala 39:24]
  reg [15:0] L0Memory_0; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_1; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_2; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_3; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_4; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_5; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_6; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_7; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_8; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_9; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_10; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_11; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_12; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_13; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_14; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_15; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_16; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_17; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_18; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_19; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_20; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_21; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_22; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_23; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_24; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_25; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_26; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_27; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_28; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_29; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_30; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_31; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_32; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_33; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_34; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_35; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_36; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_37; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_38; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_39; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_40; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_41; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_42; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_43; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_44; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_45; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_46; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_47; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_48; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_49; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_50; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_51; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_52; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_53; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_54; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_55; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_56; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_57; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_58; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_59; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_60; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_61; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_62; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_63; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_64; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_65; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_66; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_67; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_68; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_69; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_70; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_71; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_72; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_73; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_74; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_75; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_76; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_77; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_78; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_79; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_80; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_81; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_82; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_83; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_84; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_85; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_86; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_87; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_88; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_89; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_90; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_91; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_92; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_93; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_94; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_95; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_96; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_97; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_98; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_99; // @[PEArray.scala 40:21]
  reg [2:0] state; // @[PEArray.scala 100:22]
  wire  _T_3 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_12 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_16 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_22 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_31 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_41 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_342 = _T_41 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 231:12 PEArray.scala 32:8]
  wire  _GEN_349 = _T_31 ? 1'h0 : _GEN_342; // @[Conditional.scala 39:67 PEArray.scala 208:12]
  wire  _GEN_459 = _T_22 | _GEN_349; // @[Conditional.scala 39:67 PEArray.scala 32:8]
  wire  _GEN_463 = _T_16 ? 1'h0 : _GEN_459; // @[Conditional.scala 39:67]
  wire  _GEN_572 = _T_12 | _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 149:12]
  wire  sel1 = _T_3 | _GEN_572; // @[Conditional.scala 40:58 PEArray.scala 108:12]
  wire [15:0] MAC_out = FP16MAC_io_out; // @[PEArray.scala 47:21 PEArray.scala 85:11]
  wire  _GEN_465 = _T_16 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 177:12]
  wire  _GEN_580 = _T_12 | _GEN_465; // @[Conditional.scala 39:67 PEArray.scala 34:8]
  wire  sel3 = _T_3 | _GEN_580; // @[Conditional.scala 40:58 PEArray.scala 110:12]
  wire [1:0] _GEN_344 = _T_41 ? 2'h2 : 2'h0; // @[Conditional.scala 39:67 PEArray.scala 233:12 PEArray.scala 35:8]
  wire [1:0] _GEN_351 = _T_31 ? 2'h2 : _GEN_344; // @[Conditional.scala 39:67 PEArray.scala 210:12]
  wire [1:0] _GEN_461 = _T_22 ? 2'h0 : _GEN_351; // @[Conditional.scala 39:67 PEArray.scala 35:8]
  wire [1:0] _GEN_466 = _T_16 ? 2'h0 : _GEN_461; // @[Conditional.scala 39:67 PEArray.scala 178:12]
  wire [1:0] _GEN_574 = _T_12 ? 2'h1 : _GEN_466; // @[Conditional.scala 39:67]
  wire [1:0] sel4 = _T_3 ? 2'h0 : _GEN_574; // @[Conditional.scala 40:58 PEArray.scala 111:12]
  wire [15:0] _GEN_3 = sel4 == 2'h2 ? io_FromL1 : 16'h0; // @[PEArray.scala 65:28 PEArray.scala 66:15 PEArray.scala 69:15]
  wire [15:0] _GEN_4 = sel4 == 2'h1 ? io_FromAbovePE : _GEN_3; // @[PEArray.scala 62:28 PEArray.scala 63:15]
  wire [15:0] mux4out = sel4 == 2'h0 ? 16'h0 : _GEN_4; // @[PEArray.scala 59:22 PEArray.scala 60:13]
  wire [15:0] _GEN_7 = 6'h1 == L0Index ? L0Memory_1 : L0Memory_0; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_8 = 6'h2 == L0Index ? L0Memory_2 : _GEN_7; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_9 = 6'h3 == L0Index ? L0Memory_3 : _GEN_8; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_10 = 6'h4 == L0Index ? L0Memory_4 : _GEN_9; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_11 = 6'h5 == L0Index ? L0Memory_5 : _GEN_10; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_12 = 6'h6 == L0Index ? L0Memory_6 : _GEN_11; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_13 = 6'h7 == L0Index ? L0Memory_7 : _GEN_12; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_14 = 6'h8 == L0Index ? L0Memory_8 : _GEN_13; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_15 = 6'h9 == L0Index ? L0Memory_9 : _GEN_14; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_16 = 6'ha == L0Index ? L0Memory_10 : _GEN_15; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_17 = 6'hb == L0Index ? L0Memory_11 : _GEN_16; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_18 = 6'hc == L0Index ? L0Memory_12 : _GEN_17; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_19 = 6'hd == L0Index ? L0Memory_13 : _GEN_18; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_20 = 6'he == L0Index ? L0Memory_14 : _GEN_19; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_21 = 6'hf == L0Index ? L0Memory_15 : _GEN_20; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_22 = 6'h10 == L0Index ? L0Memory_16 : _GEN_21; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_23 = 6'h11 == L0Index ? L0Memory_17 : _GEN_22; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_24 = 6'h12 == L0Index ? L0Memory_18 : _GEN_23; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_25 = 6'h13 == L0Index ? L0Memory_19 : _GEN_24; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_26 = 6'h14 == L0Index ? L0Memory_20 : _GEN_25; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_27 = 6'h15 == L0Index ? L0Memory_21 : _GEN_26; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_28 = 6'h16 == L0Index ? L0Memory_22 : _GEN_27; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_29 = 6'h17 == L0Index ? L0Memory_23 : _GEN_28; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_30 = 6'h18 == L0Index ? L0Memory_24 : _GEN_29; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_31 = 6'h19 == L0Index ? L0Memory_25 : _GEN_30; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_32 = 6'h1a == L0Index ? L0Memory_26 : _GEN_31; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_33 = 6'h1b == L0Index ? L0Memory_27 : _GEN_32; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_34 = 6'h1c == L0Index ? L0Memory_28 : _GEN_33; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_35 = 6'h1d == L0Index ? L0Memory_29 : _GEN_34; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_36 = 6'h1e == L0Index ? L0Memory_30 : _GEN_35; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_37 = 6'h1f == L0Index ? L0Memory_31 : _GEN_36; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_38 = 6'h20 == L0Index ? L0Memory_32 : _GEN_37; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_39 = 6'h21 == L0Index ? L0Memory_33 : _GEN_38; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_40 = 6'h22 == L0Index ? L0Memory_34 : _GEN_39; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_41 = 6'h23 == L0Index ? L0Memory_35 : _GEN_40; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_42 = 6'h24 == L0Index ? L0Memory_36 : _GEN_41; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_43 = 6'h25 == L0Index ? L0Memory_37 : _GEN_42; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_44 = 6'h26 == L0Index ? L0Memory_38 : _GEN_43; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_45 = 6'h27 == L0Index ? L0Memory_39 : _GEN_44; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_46 = 6'h28 == L0Index ? L0Memory_40 : _GEN_45; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_47 = 6'h29 == L0Index ? L0Memory_41 : _GEN_46; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_48 = 6'h2a == L0Index ? L0Memory_42 : _GEN_47; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_49 = 6'h2b == L0Index ? L0Memory_43 : _GEN_48; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_50 = 6'h2c == L0Index ? L0Memory_44 : _GEN_49; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_51 = 6'h2d == L0Index ? L0Memory_45 : _GEN_50; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_52 = 6'h2e == L0Index ? L0Memory_46 : _GEN_51; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_53 = 6'h2f == L0Index ? L0Memory_47 : _GEN_52; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_54 = 6'h30 == L0Index ? L0Memory_48 : _GEN_53; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_55 = 6'h31 == L0Index ? L0Memory_49 : _GEN_54; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_56 = 6'h32 == L0Index ? L0Memory_50 : _GEN_55; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_57 = 6'h33 == L0Index ? L0Memory_51 : _GEN_56; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_58 = 6'h34 == L0Index ? L0Memory_52 : _GEN_57; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_59 = 6'h35 == L0Index ? L0Memory_53 : _GEN_58; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_60 = 6'h36 == L0Index ? L0Memory_54 : _GEN_59; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_61 = 6'h37 == L0Index ? L0Memory_55 : _GEN_60; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_62 = 6'h38 == L0Index ? L0Memory_56 : _GEN_61; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_63 = 6'h39 == L0Index ? L0Memory_57 : _GEN_62; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_64 = 6'h3a == L0Index ? L0Memory_58 : _GEN_63; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_65 = 6'h3b == L0Index ? L0Memory_59 : _GEN_64; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_66 = 6'h3c == L0Index ? L0Memory_60 : _GEN_65; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_67 = 6'h3d == L0Index ? L0Memory_61 : _GEN_66; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_68 = 6'h3e == L0Index ? L0Memory_62 : _GEN_67; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_69 = 6'h3f == L0Index ? L0Memory_63 : _GEN_68; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [6:0] _GEN_793 = {{1'd0}, L0Index}; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_70 = 7'h40 == _GEN_793 ? L0Memory_64 : _GEN_69; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_71 = 7'h41 == _GEN_793 ? L0Memory_65 : _GEN_70; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_72 = 7'h42 == _GEN_793 ? L0Memory_66 : _GEN_71; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_73 = 7'h43 == _GEN_793 ? L0Memory_67 : _GEN_72; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_74 = 7'h44 == _GEN_793 ? L0Memory_68 : _GEN_73; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_75 = 7'h45 == _GEN_793 ? L0Memory_69 : _GEN_74; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_76 = 7'h46 == _GEN_793 ? L0Memory_70 : _GEN_75; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_77 = 7'h47 == _GEN_793 ? L0Memory_71 : _GEN_76; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_78 = 7'h48 == _GEN_793 ? L0Memory_72 : _GEN_77; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_79 = 7'h49 == _GEN_793 ? L0Memory_73 : _GEN_78; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_80 = 7'h4a == _GEN_793 ? L0Memory_74 : _GEN_79; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_81 = 7'h4b == _GEN_793 ? L0Memory_75 : _GEN_80; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_82 = 7'h4c == _GEN_793 ? L0Memory_76 : _GEN_81; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_83 = 7'h4d == _GEN_793 ? L0Memory_77 : _GEN_82; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_84 = 7'h4e == _GEN_793 ? L0Memory_78 : _GEN_83; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_85 = 7'h4f == _GEN_793 ? L0Memory_79 : _GEN_84; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_86 = 7'h50 == _GEN_793 ? L0Memory_80 : _GEN_85; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_87 = 7'h51 == _GEN_793 ? L0Memory_81 : _GEN_86; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_88 = 7'h52 == _GEN_793 ? L0Memory_82 : _GEN_87; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_89 = 7'h53 == _GEN_793 ? L0Memory_83 : _GEN_88; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_90 = 7'h54 == _GEN_793 ? L0Memory_84 : _GEN_89; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_91 = 7'h55 == _GEN_793 ? L0Memory_85 : _GEN_90; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_92 = 7'h56 == _GEN_793 ? L0Memory_86 : _GEN_91; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_93 = 7'h57 == _GEN_793 ? L0Memory_87 : _GEN_92; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_94 = 7'h58 == _GEN_793 ? L0Memory_88 : _GEN_93; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_95 = 7'h59 == _GEN_793 ? L0Memory_89 : _GEN_94; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_96 = 7'h5a == _GEN_793 ? L0Memory_90 : _GEN_95; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_97 = 7'h5b == _GEN_793 ? L0Memory_91 : _GEN_96; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_98 = 7'h5c == _GEN_793 ? L0Memory_92 : _GEN_97; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_99 = 7'h5d == _GEN_793 ? L0Memory_93 : _GEN_98; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_100 = 7'h5e == _GEN_793 ? L0Memory_94 : _GEN_99; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_101 = 7'h5f == _GEN_793 ? L0Memory_95 : _GEN_100; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_102 = 7'h60 == _GEN_793 ? L0Memory_96 : _GEN_101; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_103 = 7'h61 == _GEN_793 ? L0Memory_97 : _GEN_102; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_104 = 7'h62 == _GEN_793 ? L0Memory_98 : _GEN_103; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_105 = 7'h63 == _GEN_793 ? L0Memory_99 : _GEN_104; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire  _GEN_575 = _T_12 ? 1'h0 : _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 157:12]
  wire  sel5 = _T_3 ? 1'h0 : _GEN_575; // @[Conditional.scala 40:58 PEArray.scala 112:12]
  reg [15:0] mux2out_reg; // @[PEArray.scala 90:28]
  reg [15:0] mux3out_reg; // @[PEArray.scala 91:28]
  reg [9:0] count; // @[PEArray.scala 101:22]
  reg [9:0] count_max; // @[PEArray.scala 102:22]
  reg [5:0] L0index_begin; // @[PEArray.scala 103:26]
  reg [5:0] GRU_out_width; // @[PEArray.scala 104:26]
  wire  _T_6 = 3'h0 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_7 = 3'h1 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_8 = 3'h2 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_9 = 3'h3 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_10 = 3'h4 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_11 = 3'h5 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_109 = _T_11 ? 3'h5 : state; // @[Conditional.scala 39:67 PEArray.scala 140:19 PEArray.scala 100:22]
  wire [2:0] _GEN_110 = _T_10 ? 3'h4 : _GEN_109; // @[Conditional.scala 39:67 PEArray.scala 136:19]
  wire [2:0] _GEN_111 = _T_9 ? 3'h3 : _GEN_110; // @[Conditional.scala 39:67 PEArray.scala 132:19]
  wire [2:0] _GEN_112 = _T_8 ? 3'h2 : _GEN_111; // @[Conditional.scala 39:67 PEArray.scala 128:19]
  wire [2:0] _GEN_113 = _T_7 ? 3'h1 : _GEN_112; // @[Conditional.scala 39:67 PEArray.scala 124:19]
  wire [7:0] _GEN_118 = io_control_signal_mask[9] ? io_control_signal_gru_out_width : {{2'd0}, GRU_out_width}; // @[PEArray.scala 116:57 PEArray.scala 145:23 PEArray.scala 104:26]
  wire [9:0] _count_T_1 = count + 10'h1; // @[PEArray.scala 162:24]
  wire [9:0] _GEN_120 = count != 10'h33 ? _count_T_1 : count; // @[PEArray.scala 161:27 PEArray.scala 162:15 PEArray.scala 101:22]
  wire [9:0] _GEN_124 = count != 10'h188 ? _count_T_1 : count; // @[PEArray.scala 183:28 PEArray.scala 184:15 PEArray.scala 101:22]
  wire [9:0] _GEN_125 = count == 10'h188 ? 10'h0 : _GEN_124; // @[PEArray.scala 186:28 PEArray.scala 187:15]
  wire [2:0] _GEN_126 = count == 10'h188 ? 3'h0 : state; // @[PEArray.scala 186:28 PEArray.scala 188:15 PEArray.scala 100:22]
  wire [9:0] _GEN_127 = count != count_max ? _count_T_1 : count; // @[PEArray.scala 192:32 PEArray.scala 193:15 PEArray.scala 101:22]
  wire [5:0] _GEN_128 = count == 10'h0 ? L0index_begin : L0Index; // @[PEArray.scala 195:26 PEArray.scala 196:17 PEArray.scala 39:24]
  wire [9:0] _T_27 = count_max - 10'h1; // @[PEArray.scala 198:51]
  wire [15:0] _GEN_129 = 6'h0 == L0Index ? io_FromL1 : L0Memory_0; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_130 = 6'h1 == L0Index ? io_FromL1 : L0Memory_1; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_131 = 6'h2 == L0Index ? io_FromL1 : L0Memory_2; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_132 = 6'h3 == L0Index ? io_FromL1 : L0Memory_3; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_133 = 6'h4 == L0Index ? io_FromL1 : L0Memory_4; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_134 = 6'h5 == L0Index ? io_FromL1 : L0Memory_5; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_135 = 6'h6 == L0Index ? io_FromL1 : L0Memory_6; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_136 = 6'h7 == L0Index ? io_FromL1 : L0Memory_7; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_137 = 6'h8 == L0Index ? io_FromL1 : L0Memory_8; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_138 = 6'h9 == L0Index ? io_FromL1 : L0Memory_9; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_139 = 6'ha == L0Index ? io_FromL1 : L0Memory_10; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_140 = 6'hb == L0Index ? io_FromL1 : L0Memory_11; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_141 = 6'hc == L0Index ? io_FromL1 : L0Memory_12; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_142 = 6'hd == L0Index ? io_FromL1 : L0Memory_13; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_143 = 6'he == L0Index ? io_FromL1 : L0Memory_14; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_144 = 6'hf == L0Index ? io_FromL1 : L0Memory_15; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_145 = 6'h10 == L0Index ? io_FromL1 : L0Memory_16; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_146 = 6'h11 == L0Index ? io_FromL1 : L0Memory_17; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_147 = 6'h12 == L0Index ? io_FromL1 : L0Memory_18; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_148 = 6'h13 == L0Index ? io_FromL1 : L0Memory_19; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_149 = 6'h14 == L0Index ? io_FromL1 : L0Memory_20; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_150 = 6'h15 == L0Index ? io_FromL1 : L0Memory_21; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_151 = 6'h16 == L0Index ? io_FromL1 : L0Memory_22; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_152 = 6'h17 == L0Index ? io_FromL1 : L0Memory_23; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_153 = 6'h18 == L0Index ? io_FromL1 : L0Memory_24; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_154 = 6'h19 == L0Index ? io_FromL1 : L0Memory_25; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_155 = 6'h1a == L0Index ? io_FromL1 : L0Memory_26; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_156 = 6'h1b == L0Index ? io_FromL1 : L0Memory_27; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_157 = 6'h1c == L0Index ? io_FromL1 : L0Memory_28; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_158 = 6'h1d == L0Index ? io_FromL1 : L0Memory_29; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_159 = 6'h1e == L0Index ? io_FromL1 : L0Memory_30; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_160 = 6'h1f == L0Index ? io_FromL1 : L0Memory_31; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_161 = 6'h20 == L0Index ? io_FromL1 : L0Memory_32; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_162 = 6'h21 == L0Index ? io_FromL1 : L0Memory_33; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_163 = 6'h22 == L0Index ? io_FromL1 : L0Memory_34; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_164 = 6'h23 == L0Index ? io_FromL1 : L0Memory_35; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_165 = 6'h24 == L0Index ? io_FromL1 : L0Memory_36; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_166 = 6'h25 == L0Index ? io_FromL1 : L0Memory_37; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_167 = 6'h26 == L0Index ? io_FromL1 : L0Memory_38; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_168 = 6'h27 == L0Index ? io_FromL1 : L0Memory_39; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_169 = 6'h28 == L0Index ? io_FromL1 : L0Memory_40; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_170 = 6'h29 == L0Index ? io_FromL1 : L0Memory_41; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_171 = 6'h2a == L0Index ? io_FromL1 : L0Memory_42; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_172 = 6'h2b == L0Index ? io_FromL1 : L0Memory_43; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_173 = 6'h2c == L0Index ? io_FromL1 : L0Memory_44; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_174 = 6'h2d == L0Index ? io_FromL1 : L0Memory_45; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_175 = 6'h2e == L0Index ? io_FromL1 : L0Memory_46; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_176 = 6'h2f == L0Index ? io_FromL1 : L0Memory_47; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_177 = 6'h30 == L0Index ? io_FromL1 : L0Memory_48; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_178 = 6'h31 == L0Index ? io_FromL1 : L0Memory_49; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_179 = 6'h32 == L0Index ? io_FromL1 : L0Memory_50; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_180 = 6'h33 == L0Index ? io_FromL1 : L0Memory_51; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_181 = 6'h34 == L0Index ? io_FromL1 : L0Memory_52; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_182 = 6'h35 == L0Index ? io_FromL1 : L0Memory_53; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_183 = 6'h36 == L0Index ? io_FromL1 : L0Memory_54; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_184 = 6'h37 == L0Index ? io_FromL1 : L0Memory_55; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_185 = 6'h38 == L0Index ? io_FromL1 : L0Memory_56; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_186 = 6'h39 == L0Index ? io_FromL1 : L0Memory_57; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_187 = 6'h3a == L0Index ? io_FromL1 : L0Memory_58; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_188 = 6'h3b == L0Index ? io_FromL1 : L0Memory_59; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_189 = 6'h3c == L0Index ? io_FromL1 : L0Memory_60; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_190 = 6'h3d == L0Index ? io_FromL1 : L0Memory_61; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_191 = 6'h3e == L0Index ? io_FromL1 : L0Memory_62; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_192 = 6'h3f == L0Index ? io_FromL1 : L0Memory_63; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_193 = 7'h40 == _GEN_793 ? io_FromL1 : L0Memory_64; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_194 = 7'h41 == _GEN_793 ? io_FromL1 : L0Memory_65; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_195 = 7'h42 == _GEN_793 ? io_FromL1 : L0Memory_66; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_196 = 7'h43 == _GEN_793 ? io_FromL1 : L0Memory_67; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_197 = 7'h44 == _GEN_793 ? io_FromL1 : L0Memory_68; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_198 = 7'h45 == _GEN_793 ? io_FromL1 : L0Memory_69; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_199 = 7'h46 == _GEN_793 ? io_FromL1 : L0Memory_70; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_200 = 7'h47 == _GEN_793 ? io_FromL1 : L0Memory_71; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_201 = 7'h48 == _GEN_793 ? io_FromL1 : L0Memory_72; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_202 = 7'h49 == _GEN_793 ? io_FromL1 : L0Memory_73; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_203 = 7'h4a == _GEN_793 ? io_FromL1 : L0Memory_74; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_204 = 7'h4b == _GEN_793 ? io_FromL1 : L0Memory_75; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_205 = 7'h4c == _GEN_793 ? io_FromL1 : L0Memory_76; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_206 = 7'h4d == _GEN_793 ? io_FromL1 : L0Memory_77; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_207 = 7'h4e == _GEN_793 ? io_FromL1 : L0Memory_78; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_208 = 7'h4f == _GEN_793 ? io_FromL1 : L0Memory_79; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_209 = 7'h50 == _GEN_793 ? io_FromL1 : L0Memory_80; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_210 = 7'h51 == _GEN_793 ? io_FromL1 : L0Memory_81; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_211 = 7'h52 == _GEN_793 ? io_FromL1 : L0Memory_82; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_212 = 7'h53 == _GEN_793 ? io_FromL1 : L0Memory_83; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_213 = 7'h54 == _GEN_793 ? io_FromL1 : L0Memory_84; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_214 = 7'h55 == _GEN_793 ? io_FromL1 : L0Memory_85; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_215 = 7'h56 == _GEN_793 ? io_FromL1 : L0Memory_86; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_216 = 7'h57 == _GEN_793 ? io_FromL1 : L0Memory_87; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_217 = 7'h58 == _GEN_793 ? io_FromL1 : L0Memory_88; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_218 = 7'h59 == _GEN_793 ? io_FromL1 : L0Memory_89; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_219 = 7'h5a == _GEN_793 ? io_FromL1 : L0Memory_90; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_220 = 7'h5b == _GEN_793 ? io_FromL1 : L0Memory_91; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_221 = 7'h5c == _GEN_793 ? io_FromL1 : L0Memory_92; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_222 = 7'h5d == _GEN_793 ? io_FromL1 : L0Memory_93; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_223 = 7'h5e == _GEN_793 ? io_FromL1 : L0Memory_94; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_224 = 7'h5f == _GEN_793 ? io_FromL1 : L0Memory_95; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_225 = 7'h60 == _GEN_793 ? io_FromL1 : L0Memory_96; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_226 = 7'h61 == _GEN_793 ? io_FromL1 : L0Memory_97; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_227 = 7'h62 == _GEN_793 ? io_FromL1 : L0Memory_98; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_228 = 7'h63 == _GEN_793 ? io_FromL1 : L0Memory_99; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [5:0] _L0Index_T_2 = L0Index + 6'h1; // @[PEArray.scala 200:28]
  wire [15:0] _GEN_229 = count >= 10'h1 & count <= _T_27 ? _GEN_129 : L0Memory_0; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_230 = count >= 10'h1 & count <= _T_27 ? _GEN_130 : L0Memory_1; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_231 = count >= 10'h1 & count <= _T_27 ? _GEN_131 : L0Memory_2; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_232 = count >= 10'h1 & count <= _T_27 ? _GEN_132 : L0Memory_3; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_233 = count >= 10'h1 & count <= _T_27 ? _GEN_133 : L0Memory_4; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_234 = count >= 10'h1 & count <= _T_27 ? _GEN_134 : L0Memory_5; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_235 = count >= 10'h1 & count <= _T_27 ? _GEN_135 : L0Memory_6; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_236 = count >= 10'h1 & count <= _T_27 ? _GEN_136 : L0Memory_7; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_237 = count >= 10'h1 & count <= _T_27 ? _GEN_137 : L0Memory_8; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_238 = count >= 10'h1 & count <= _T_27 ? _GEN_138 : L0Memory_9; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_239 = count >= 10'h1 & count <= _T_27 ? _GEN_139 : L0Memory_10; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_240 = count >= 10'h1 & count <= _T_27 ? _GEN_140 : L0Memory_11; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_241 = count >= 10'h1 & count <= _T_27 ? _GEN_141 : L0Memory_12; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_242 = count >= 10'h1 & count <= _T_27 ? _GEN_142 : L0Memory_13; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_243 = count >= 10'h1 & count <= _T_27 ? _GEN_143 : L0Memory_14; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_244 = count >= 10'h1 & count <= _T_27 ? _GEN_144 : L0Memory_15; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_245 = count >= 10'h1 & count <= _T_27 ? _GEN_145 : L0Memory_16; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_246 = count >= 10'h1 & count <= _T_27 ? _GEN_146 : L0Memory_17; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_247 = count >= 10'h1 & count <= _T_27 ? _GEN_147 : L0Memory_18; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_248 = count >= 10'h1 & count <= _T_27 ? _GEN_148 : L0Memory_19; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_249 = count >= 10'h1 & count <= _T_27 ? _GEN_149 : L0Memory_20; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_250 = count >= 10'h1 & count <= _T_27 ? _GEN_150 : L0Memory_21; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_251 = count >= 10'h1 & count <= _T_27 ? _GEN_151 : L0Memory_22; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_252 = count >= 10'h1 & count <= _T_27 ? _GEN_152 : L0Memory_23; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_253 = count >= 10'h1 & count <= _T_27 ? _GEN_153 : L0Memory_24; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_254 = count >= 10'h1 & count <= _T_27 ? _GEN_154 : L0Memory_25; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_255 = count >= 10'h1 & count <= _T_27 ? _GEN_155 : L0Memory_26; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_256 = count >= 10'h1 & count <= _T_27 ? _GEN_156 : L0Memory_27; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_257 = count >= 10'h1 & count <= _T_27 ? _GEN_157 : L0Memory_28; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_258 = count >= 10'h1 & count <= _T_27 ? _GEN_158 : L0Memory_29; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_259 = count >= 10'h1 & count <= _T_27 ? _GEN_159 : L0Memory_30; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_260 = count >= 10'h1 & count <= _T_27 ? _GEN_160 : L0Memory_31; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_261 = count >= 10'h1 & count <= _T_27 ? _GEN_161 : L0Memory_32; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_262 = count >= 10'h1 & count <= _T_27 ? _GEN_162 : L0Memory_33; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_263 = count >= 10'h1 & count <= _T_27 ? _GEN_163 : L0Memory_34; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_264 = count >= 10'h1 & count <= _T_27 ? _GEN_164 : L0Memory_35; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_265 = count >= 10'h1 & count <= _T_27 ? _GEN_165 : L0Memory_36; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_266 = count >= 10'h1 & count <= _T_27 ? _GEN_166 : L0Memory_37; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_267 = count >= 10'h1 & count <= _T_27 ? _GEN_167 : L0Memory_38; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_268 = count >= 10'h1 & count <= _T_27 ? _GEN_168 : L0Memory_39; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_269 = count >= 10'h1 & count <= _T_27 ? _GEN_169 : L0Memory_40; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_270 = count >= 10'h1 & count <= _T_27 ? _GEN_170 : L0Memory_41; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_271 = count >= 10'h1 & count <= _T_27 ? _GEN_171 : L0Memory_42; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_272 = count >= 10'h1 & count <= _T_27 ? _GEN_172 : L0Memory_43; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_273 = count >= 10'h1 & count <= _T_27 ? _GEN_173 : L0Memory_44; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_274 = count >= 10'h1 & count <= _T_27 ? _GEN_174 : L0Memory_45; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_275 = count >= 10'h1 & count <= _T_27 ? _GEN_175 : L0Memory_46; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_276 = count >= 10'h1 & count <= _T_27 ? _GEN_176 : L0Memory_47; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_277 = count >= 10'h1 & count <= _T_27 ? _GEN_177 : L0Memory_48; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_278 = count >= 10'h1 & count <= _T_27 ? _GEN_178 : L0Memory_49; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_279 = count >= 10'h1 & count <= _T_27 ? _GEN_179 : L0Memory_50; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_280 = count >= 10'h1 & count <= _T_27 ? _GEN_180 : L0Memory_51; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_281 = count >= 10'h1 & count <= _T_27 ? _GEN_181 : L0Memory_52; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_282 = count >= 10'h1 & count <= _T_27 ? _GEN_182 : L0Memory_53; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_283 = count >= 10'h1 & count <= _T_27 ? _GEN_183 : L0Memory_54; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_284 = count >= 10'h1 & count <= _T_27 ? _GEN_184 : L0Memory_55; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_285 = count >= 10'h1 & count <= _T_27 ? _GEN_185 : L0Memory_56; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_286 = count >= 10'h1 & count <= _T_27 ? _GEN_186 : L0Memory_57; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_287 = count >= 10'h1 & count <= _T_27 ? _GEN_187 : L0Memory_58; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_288 = count >= 10'h1 & count <= _T_27 ? _GEN_188 : L0Memory_59; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_289 = count >= 10'h1 & count <= _T_27 ? _GEN_189 : L0Memory_60; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_290 = count >= 10'h1 & count <= _T_27 ? _GEN_190 : L0Memory_61; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_291 = count >= 10'h1 & count <= _T_27 ? _GEN_191 : L0Memory_62; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_292 = count >= 10'h1 & count <= _T_27 ? _GEN_192 : L0Memory_63; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_293 = count >= 10'h1 & count <= _T_27 ? _GEN_193 : L0Memory_64; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_294 = count >= 10'h1 & count <= _T_27 ? _GEN_194 : L0Memory_65; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_295 = count >= 10'h1 & count <= _T_27 ? _GEN_195 : L0Memory_66; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_296 = count >= 10'h1 & count <= _T_27 ? _GEN_196 : L0Memory_67; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_297 = count >= 10'h1 & count <= _T_27 ? _GEN_197 : L0Memory_68; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_298 = count >= 10'h1 & count <= _T_27 ? _GEN_198 : L0Memory_69; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_299 = count >= 10'h1 & count <= _T_27 ? _GEN_199 : L0Memory_70; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_300 = count >= 10'h1 & count <= _T_27 ? _GEN_200 : L0Memory_71; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_301 = count >= 10'h1 & count <= _T_27 ? _GEN_201 : L0Memory_72; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_302 = count >= 10'h1 & count <= _T_27 ? _GEN_202 : L0Memory_73; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_303 = count >= 10'h1 & count <= _T_27 ? _GEN_203 : L0Memory_74; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_304 = count >= 10'h1 & count <= _T_27 ? _GEN_204 : L0Memory_75; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_305 = count >= 10'h1 & count <= _T_27 ? _GEN_205 : L0Memory_76; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_306 = count >= 10'h1 & count <= _T_27 ? _GEN_206 : L0Memory_77; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_307 = count >= 10'h1 & count <= _T_27 ? _GEN_207 : L0Memory_78; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_308 = count >= 10'h1 & count <= _T_27 ? _GEN_208 : L0Memory_79; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_309 = count >= 10'h1 & count <= _T_27 ? _GEN_209 : L0Memory_80; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_310 = count >= 10'h1 & count <= _T_27 ? _GEN_210 : L0Memory_81; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_311 = count >= 10'h1 & count <= _T_27 ? _GEN_211 : L0Memory_82; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_312 = count >= 10'h1 & count <= _T_27 ? _GEN_212 : L0Memory_83; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_313 = count >= 10'h1 & count <= _T_27 ? _GEN_213 : L0Memory_84; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_314 = count >= 10'h1 & count <= _T_27 ? _GEN_214 : L0Memory_85; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_315 = count >= 10'h1 & count <= _T_27 ? _GEN_215 : L0Memory_86; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_316 = count >= 10'h1 & count <= _T_27 ? _GEN_216 : L0Memory_87; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_317 = count >= 10'h1 & count <= _T_27 ? _GEN_217 : L0Memory_88; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_318 = count >= 10'h1 & count <= _T_27 ? _GEN_218 : L0Memory_89; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_319 = count >= 10'h1 & count <= _T_27 ? _GEN_219 : L0Memory_90; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_320 = count >= 10'h1 & count <= _T_27 ? _GEN_220 : L0Memory_91; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_321 = count >= 10'h1 & count <= _T_27 ? _GEN_221 : L0Memory_92; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_322 = count >= 10'h1 & count <= _T_27 ? _GEN_222 : L0Memory_93; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_323 = count >= 10'h1 & count <= _T_27 ? _GEN_223 : L0Memory_94; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_324 = count >= 10'h1 & count <= _T_27 ? _GEN_224 : L0Memory_95; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_325 = count >= 10'h1 & count <= _T_27 ? _GEN_225 : L0Memory_96; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_326 = count >= 10'h1 & count <= _T_27 ? _GEN_226 : L0Memory_97; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_327 = count >= 10'h1 & count <= _T_27 ? _GEN_227 : L0Memory_98; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_328 = count >= 10'h1 & count <= _T_27 ? _GEN_228 : L0Memory_99; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [5:0] _GEN_329 = count >= 10'h1 & count <= _T_27 ? _L0Index_T_2 : _GEN_128; // @[PEArray.scala 198:59 PEArray.scala 200:17]
  wire [9:0] _GEN_330 = count == count_max ? 10'h0 : _GEN_127; // @[PEArray.scala 202:32 PEArray.scala 203:15]
  wire [2:0] _GEN_331 = count == count_max ? 3'h0 : state; // @[PEArray.scala 202:32 PEArray.scala 204:15 PEArray.scala 100:22]
  wire [9:0] _GEN_865 = {{4'd0}, GRU_out_width}; // @[PEArray.scala 220:19]
  wire [9:0] _GEN_0 = count % _GEN_865; // @[PEArray.scala 220:19]
  wire [5:0] _T_36 = _GEN_0[5:0]; // @[PEArray.scala 220:19]
  wire [5:0] _T_38 = GRU_out_width - 6'h1; // @[PEArray.scala 220:55]
  wire [5:0] _GEN_334 = _T_36 == _T_38 ? _L0Index_T_2 : L0index_begin; // @[PEArray.scala 220:62 PEArray.scala 221:17 PEArray.scala 214:15]
  wire [5:0] _GEN_346 = _T_41 ? _GEN_334 : L0Index; // @[Conditional.scala 39:67 PEArray.scala 39:24]
  wire [9:0] _GEN_347 = _T_41 ? _GEN_330 : count; // @[Conditional.scala 39:67 PEArray.scala 101:22]
  wire [2:0] _GEN_348 = _T_41 ? _GEN_331 : state; // @[Conditional.scala 39:67 PEArray.scala 100:22]
  wire [5:0] _GEN_353 = _T_31 ? _GEN_334 : _GEN_346; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_354 = _T_31 ? _GEN_330 : _GEN_347; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_355 = _T_31 ? _GEN_331 : _GEN_348; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_356 = _T_22 ? _GEN_330 : _GEN_354; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_357 = _T_22 ? _GEN_329 : _GEN_353; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_458 = _T_22 ? _GEN_331 : _GEN_355; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_690 = _T_3 ? _GEN_118 : {{2'd0}, GRU_out_width}; // @[Conditional.scala 40:58 PEArray.scala 104:26]
  FP16MulAdder FP16MAC ( // @[PEArray.scala 72:23]
    .io_a(FP16MAC_io_a),
    .io_b(FP16MAC_io_b),
    .io_c(FP16MAC_io_c),
    .io_out(FP16MAC_io_out)
  );
  assign io_ToRightPE = mux3out_reg; // @[PEArray.scala 95:16]
  assign io_ToBelowPE = mux2out_reg; // @[PEArray.scala 94:16]
  assign FP16MAC_io_a = sel1 ? io_FromL1 : io_FromLeftPE; // @[PEArray.scala 50:14 PEArray.scala 50:23 PEArray.scala 51:24]
  assign FP16MAC_io_b = sel5 ? mux4out : _GEN_105; // @[PEArray.scala 77:13 PEArray.scala 78:18 PEArray.scala 81:18]
  assign FP16MAC_io_c = sel5 ? _GEN_105 : mux4out; // @[PEArray.scala 77:13 PEArray.scala 79:18 PEArray.scala 82:18]
  always @(posedge clock) begin
    if (reset) begin // @[PEArray.scala 39:24]
      L0Index <= 6'h0; // @[PEArray.scala 39:24]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h2; // @[PEArray.scala 159:15]
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h5; // @[PEArray.scala 181:15]
      end else begin
        L0Index <= _GEN_357;
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_0 <= _GEN_229;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_1 <= _GEN_230;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_2 <= _GEN_231;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_3 <= _GEN_232;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_4 <= _GEN_233;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_5 <= _GEN_234;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_6 <= _GEN_235;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_7 <= _GEN_236;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_8 <= _GEN_237;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_9 <= _GEN_238;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_10 <= _GEN_239;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_11 <= _GEN_240;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_12 <= _GEN_241;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_13 <= _GEN_242;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_14 <= _GEN_243;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_15 <= _GEN_244;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_16 <= _GEN_245;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_17 <= _GEN_246;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_18 <= _GEN_247;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_19 <= _GEN_248;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_20 <= _GEN_249;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_21 <= _GEN_250;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_22 <= _GEN_251;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_23 <= _GEN_252;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_24 <= _GEN_253;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_25 <= _GEN_254;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_26 <= _GEN_255;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_27 <= _GEN_256;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_28 <= _GEN_257;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_29 <= _GEN_258;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_30 <= _GEN_259;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_31 <= _GEN_260;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_32 <= _GEN_261;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_33 <= _GEN_262;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_34 <= _GEN_263;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_35 <= _GEN_264;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_36 <= _GEN_265;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_37 <= _GEN_266;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_38 <= _GEN_267;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_39 <= _GEN_268;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_40 <= _GEN_269;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_41 <= _GEN_270;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_42 <= _GEN_271;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_43 <= _GEN_272;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_44 <= _GEN_273;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_45 <= _GEN_274;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_46 <= _GEN_275;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_47 <= _GEN_276;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_48 <= _GEN_277;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_49 <= _GEN_278;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_50 <= _GEN_279;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_51 <= _GEN_280;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_52 <= _GEN_281;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_53 <= _GEN_282;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_54 <= _GEN_283;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_55 <= _GEN_284;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_56 <= _GEN_285;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_57 <= _GEN_286;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_58 <= _GEN_287;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_59 <= _GEN_288;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_60 <= _GEN_289;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_61 <= _GEN_290;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_62 <= _GEN_291;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_63 <= _GEN_292;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_64 <= _GEN_293;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_65 <= _GEN_294;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_66 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_67 <= _GEN_296;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_68 <= _GEN_297;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_69 <= _GEN_298;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_70 <= _GEN_299;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_71 <= _GEN_300;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_72 <= _GEN_301;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_73 <= _GEN_302;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_74 <= _GEN_303;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_75 <= _GEN_304;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_76 <= _GEN_305;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_77 <= _GEN_306;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_78 <= _GEN_307;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_79 <= _GEN_308;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_80 <= _GEN_309;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_81 <= _GEN_310;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_82 <= _GEN_311;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_83 <= _GEN_312;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_84 <= _GEN_313;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_85 <= _GEN_314;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_86 <= _GEN_315;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_87 <= _GEN_316;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_88 <= _GEN_317;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_89 <= _GEN_318;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_90 <= _GEN_319;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_91 <= _GEN_320;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_92 <= _GEN_321;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_93 <= _GEN_322;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_94 <= _GEN_323;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_95 <= _GEN_324;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_96 <= _GEN_325;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_97 <= _GEN_326;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_98 <= _GEN_327;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_99 <= _GEN_328;
          end
        end
      end
    end
    if (reset) begin // @[PEArray.scala 100:22]
      state <= 3'h0; // @[PEArray.scala 100:22]
    end else if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[9]) begin // @[PEArray.scala 116:57]
        if (_T_6) begin // @[Conditional.scala 40:58]
          state <= 3'h0; // @[PEArray.scala 120:19]
        end else begin
          state <= _GEN_113;
        end
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      if (count == 10'h33) begin // @[PEArray.scala 164:27]
        state <= 3'h0; // @[PEArray.scala 166:15]
      end
    end else if (_T_16) begin // @[Conditional.scala 39:67]
      state <= _GEN_126;
    end else begin
      state <= _GEN_458;
    end
    if (reset) begin // @[PEArray.scala 90:28]
      mux2out_reg <= 16'h0; // @[PEArray.scala 90:28]
    end else begin
      mux2out_reg <= MAC_out; // @[PEArray.scala 90:28]
    end
    if (reset) begin // @[PEArray.scala 91:28]
      mux3out_reg <= 16'h0; // @[PEArray.scala 91:28]
    end else if (sel3) begin // @[PEArray.scala 56:14]
      mux3out_reg <= MAC_out; // @[PEArray.scala 56:23]
    end else if (sel1) begin // @[PEArray.scala 50:14]
      mux3out_reg <= io_FromL1; // @[PEArray.scala 50:23]
    end else begin
      mux3out_reg <= io_FromLeftPE; // @[PEArray.scala 51:24]
    end
    if (reset) begin // @[PEArray.scala 101:22]
      count <= 10'h0; // @[PEArray.scala 101:22]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        if (count == 10'h33) begin // @[PEArray.scala 164:27]
          count <= 10'h0; // @[PEArray.scala 165:15]
        end else begin
          count <= _GEN_120;
        end
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        count <= _GEN_125;
      end else begin
        count <= _GEN_356;
      end
    end
    if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[9]) begin // @[PEArray.scala 116:57]
        count_max <= io_control_signal_count; // @[PEArray.scala 143:19]
      end
    end
    if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[9]) begin // @[PEArray.scala 116:57]
        L0index_begin <= io_control_signal_L0index; // @[PEArray.scala 144:23]
      end
    end
    GRU_out_width <= _GEN_690[5:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  L0Index = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  L0Memory_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  L0Memory_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  L0Memory_2 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  L0Memory_3 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  L0Memory_4 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  L0Memory_5 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  L0Memory_6 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  L0Memory_7 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  L0Memory_8 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  L0Memory_9 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  L0Memory_10 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  L0Memory_11 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  L0Memory_12 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  L0Memory_13 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  L0Memory_14 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  L0Memory_15 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  L0Memory_16 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  L0Memory_17 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  L0Memory_18 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  L0Memory_19 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  L0Memory_20 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  L0Memory_21 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  L0Memory_22 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  L0Memory_23 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  L0Memory_24 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  L0Memory_25 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  L0Memory_26 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  L0Memory_27 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  L0Memory_28 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  L0Memory_29 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  L0Memory_30 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  L0Memory_31 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  L0Memory_32 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  L0Memory_33 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  L0Memory_34 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  L0Memory_35 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  L0Memory_36 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  L0Memory_37 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  L0Memory_38 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  L0Memory_39 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  L0Memory_40 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  L0Memory_41 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  L0Memory_42 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  L0Memory_43 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  L0Memory_44 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  L0Memory_45 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  L0Memory_46 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  L0Memory_47 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  L0Memory_48 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  L0Memory_49 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  L0Memory_50 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  L0Memory_51 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  L0Memory_52 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  L0Memory_53 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  L0Memory_54 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  L0Memory_55 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  L0Memory_56 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  L0Memory_57 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  L0Memory_58 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  L0Memory_59 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  L0Memory_60 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  L0Memory_61 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  L0Memory_62 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  L0Memory_63 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  L0Memory_64 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  L0Memory_65 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  L0Memory_66 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  L0Memory_67 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  L0Memory_68 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  L0Memory_69 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  L0Memory_70 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  L0Memory_71 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  L0Memory_72 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  L0Memory_73 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  L0Memory_74 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  L0Memory_75 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  L0Memory_76 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  L0Memory_77 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  L0Memory_78 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  L0Memory_79 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  L0Memory_80 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  L0Memory_81 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  L0Memory_82 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  L0Memory_83 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  L0Memory_84 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  L0Memory_85 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  L0Memory_86 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  L0Memory_87 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  L0Memory_88 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  L0Memory_89 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  L0Memory_90 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  L0Memory_91 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  L0Memory_92 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  L0Memory_93 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  L0Memory_94 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  L0Memory_95 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  L0Memory_96 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  L0Memory_97 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  L0Memory_98 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  L0Memory_99 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  state = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  mux2out_reg = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  mux3out_reg = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  count = _RAND_104[9:0];
  _RAND_105 = {1{`RANDOM}};
  count_max = _RAND_105[9:0];
  _RAND_106 = {1{`RANDOM}};
  L0index_begin = _RAND_106[5:0];
  _RAND_107 = {1{`RANDOM}};
  GRU_out_width = _RAND_107[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PE_9(
  input         clock,
  input         reset,
  input  [15:0] io_FromAbovePE,
  input  [15:0] io_FromLeftPE,
  input  [15:0] io_FromL1,
  input  [11:0] io_control_signal_mask,
  output [15:0] io_ToRightPE,
  output [15:0] io_ToBelowPE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] FP16MAC_io_a; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_b; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_c; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_out; // @[PEArray.scala 72:23]
  reg [5:0] L0Index; // @[PEArray.scala 39:24]
  reg [15:0] L0Memory_0; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_1; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_2; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_3; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_4; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_5; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_6; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_7; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_8; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_9; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_10; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_11; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_12; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_13; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_14; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_15; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_16; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_17; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_18; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_19; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_20; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_21; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_22; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_23; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_24; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_25; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_26; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_27; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_28; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_29; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_30; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_31; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_32; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_33; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_34; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_35; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_36; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_37; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_38; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_39; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_40; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_41; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_42; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_43; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_44; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_45; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_46; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_47; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_48; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_49; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_50; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_51; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_52; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_53; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_54; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_55; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_56; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_57; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_58; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_59; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_60; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_61; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_62; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_63; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_64; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_65; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_66; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_67; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_68; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_69; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_70; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_71; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_72; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_73; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_74; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_75; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_76; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_77; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_78; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_79; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_80; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_81; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_82; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_83; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_84; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_85; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_86; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_87; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_88; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_89; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_90; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_91; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_92; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_93; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_94; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_95; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_96; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_97; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_98; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_99; // @[PEArray.scala 40:21]
  reg [2:0] state; // @[PEArray.scala 100:22]
  wire  _T_3 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_12 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_16 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_22 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_31 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_41 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_342 = _T_41 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 231:12 PEArray.scala 32:8]
  wire  _GEN_349 = _T_31 ? 1'h0 : _GEN_342; // @[Conditional.scala 39:67 PEArray.scala 208:12]
  wire  _GEN_459 = _T_22 | _GEN_349; // @[Conditional.scala 39:67 PEArray.scala 32:8]
  wire  _GEN_463 = _T_16 ? 1'h0 : _GEN_459; // @[Conditional.scala 39:67]
  wire  _GEN_572 = _T_12 | _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 149:12]
  wire  sel1 = _T_3 | _GEN_572; // @[Conditional.scala 40:58 PEArray.scala 108:12]
  wire [15:0] MAC_out = FP16MAC_io_out; // @[PEArray.scala 47:21 PEArray.scala 85:11]
  wire  _GEN_465 = _T_16 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 177:12]
  wire  _GEN_580 = _T_12 | _GEN_465; // @[Conditional.scala 39:67 PEArray.scala 34:8]
  wire  sel3 = _T_3 | _GEN_580; // @[Conditional.scala 40:58 PEArray.scala 110:12]
  wire [1:0] _GEN_344 = _T_41 ? 2'h2 : 2'h0; // @[Conditional.scala 39:67 PEArray.scala 233:12 PEArray.scala 35:8]
  wire [1:0] _GEN_351 = _T_31 ? 2'h2 : _GEN_344; // @[Conditional.scala 39:67 PEArray.scala 210:12]
  wire [1:0] _GEN_461 = _T_22 ? 2'h0 : _GEN_351; // @[Conditional.scala 39:67 PEArray.scala 35:8]
  wire [1:0] _GEN_466 = _T_16 ? 2'h0 : _GEN_461; // @[Conditional.scala 39:67 PEArray.scala 178:12]
  wire [1:0] _GEN_574 = _T_12 ? 2'h0 : _GEN_466; // @[Conditional.scala 39:67]
  wire [1:0] sel4 = _T_3 ? 2'h0 : _GEN_574; // @[Conditional.scala 40:58 PEArray.scala 111:12]
  wire [15:0] _GEN_3 = sel4 == 2'h2 ? io_FromL1 : 16'h0; // @[PEArray.scala 65:28 PEArray.scala 66:15 PEArray.scala 69:15]
  wire [15:0] _GEN_4 = sel4 == 2'h1 ? io_FromAbovePE : _GEN_3; // @[PEArray.scala 62:28 PEArray.scala 63:15]
  wire [15:0] mux4out = sel4 == 2'h0 ? 16'h0 : _GEN_4; // @[PEArray.scala 59:22 PEArray.scala 60:13]
  wire [15:0] _GEN_7 = 6'h1 == L0Index ? L0Memory_1 : L0Memory_0; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_8 = 6'h2 == L0Index ? L0Memory_2 : _GEN_7; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_9 = 6'h3 == L0Index ? L0Memory_3 : _GEN_8; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_10 = 6'h4 == L0Index ? L0Memory_4 : _GEN_9; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_11 = 6'h5 == L0Index ? L0Memory_5 : _GEN_10; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_12 = 6'h6 == L0Index ? L0Memory_6 : _GEN_11; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_13 = 6'h7 == L0Index ? L0Memory_7 : _GEN_12; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_14 = 6'h8 == L0Index ? L0Memory_8 : _GEN_13; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_15 = 6'h9 == L0Index ? L0Memory_9 : _GEN_14; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_16 = 6'ha == L0Index ? L0Memory_10 : _GEN_15; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_17 = 6'hb == L0Index ? L0Memory_11 : _GEN_16; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_18 = 6'hc == L0Index ? L0Memory_12 : _GEN_17; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_19 = 6'hd == L0Index ? L0Memory_13 : _GEN_18; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_20 = 6'he == L0Index ? L0Memory_14 : _GEN_19; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_21 = 6'hf == L0Index ? L0Memory_15 : _GEN_20; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_22 = 6'h10 == L0Index ? L0Memory_16 : _GEN_21; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_23 = 6'h11 == L0Index ? L0Memory_17 : _GEN_22; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_24 = 6'h12 == L0Index ? L0Memory_18 : _GEN_23; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_25 = 6'h13 == L0Index ? L0Memory_19 : _GEN_24; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_26 = 6'h14 == L0Index ? L0Memory_20 : _GEN_25; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_27 = 6'h15 == L0Index ? L0Memory_21 : _GEN_26; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_28 = 6'h16 == L0Index ? L0Memory_22 : _GEN_27; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_29 = 6'h17 == L0Index ? L0Memory_23 : _GEN_28; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_30 = 6'h18 == L0Index ? L0Memory_24 : _GEN_29; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_31 = 6'h19 == L0Index ? L0Memory_25 : _GEN_30; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_32 = 6'h1a == L0Index ? L0Memory_26 : _GEN_31; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_33 = 6'h1b == L0Index ? L0Memory_27 : _GEN_32; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_34 = 6'h1c == L0Index ? L0Memory_28 : _GEN_33; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_35 = 6'h1d == L0Index ? L0Memory_29 : _GEN_34; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_36 = 6'h1e == L0Index ? L0Memory_30 : _GEN_35; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_37 = 6'h1f == L0Index ? L0Memory_31 : _GEN_36; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_38 = 6'h20 == L0Index ? L0Memory_32 : _GEN_37; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_39 = 6'h21 == L0Index ? L0Memory_33 : _GEN_38; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_40 = 6'h22 == L0Index ? L0Memory_34 : _GEN_39; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_41 = 6'h23 == L0Index ? L0Memory_35 : _GEN_40; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_42 = 6'h24 == L0Index ? L0Memory_36 : _GEN_41; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_43 = 6'h25 == L0Index ? L0Memory_37 : _GEN_42; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_44 = 6'h26 == L0Index ? L0Memory_38 : _GEN_43; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_45 = 6'h27 == L0Index ? L0Memory_39 : _GEN_44; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_46 = 6'h28 == L0Index ? L0Memory_40 : _GEN_45; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_47 = 6'h29 == L0Index ? L0Memory_41 : _GEN_46; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_48 = 6'h2a == L0Index ? L0Memory_42 : _GEN_47; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_49 = 6'h2b == L0Index ? L0Memory_43 : _GEN_48; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_50 = 6'h2c == L0Index ? L0Memory_44 : _GEN_49; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_51 = 6'h2d == L0Index ? L0Memory_45 : _GEN_50; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_52 = 6'h2e == L0Index ? L0Memory_46 : _GEN_51; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_53 = 6'h2f == L0Index ? L0Memory_47 : _GEN_52; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_54 = 6'h30 == L0Index ? L0Memory_48 : _GEN_53; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_55 = 6'h31 == L0Index ? L0Memory_49 : _GEN_54; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_56 = 6'h32 == L0Index ? L0Memory_50 : _GEN_55; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_57 = 6'h33 == L0Index ? L0Memory_51 : _GEN_56; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_58 = 6'h34 == L0Index ? L0Memory_52 : _GEN_57; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_59 = 6'h35 == L0Index ? L0Memory_53 : _GEN_58; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_60 = 6'h36 == L0Index ? L0Memory_54 : _GEN_59; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_61 = 6'h37 == L0Index ? L0Memory_55 : _GEN_60; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_62 = 6'h38 == L0Index ? L0Memory_56 : _GEN_61; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_63 = 6'h39 == L0Index ? L0Memory_57 : _GEN_62; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_64 = 6'h3a == L0Index ? L0Memory_58 : _GEN_63; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_65 = 6'h3b == L0Index ? L0Memory_59 : _GEN_64; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_66 = 6'h3c == L0Index ? L0Memory_60 : _GEN_65; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_67 = 6'h3d == L0Index ? L0Memory_61 : _GEN_66; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_68 = 6'h3e == L0Index ? L0Memory_62 : _GEN_67; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_69 = 6'h3f == L0Index ? L0Memory_63 : _GEN_68; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [6:0] _GEN_793 = {{1'd0}, L0Index}; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_70 = 7'h40 == _GEN_793 ? L0Memory_64 : _GEN_69; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_71 = 7'h41 == _GEN_793 ? L0Memory_65 : _GEN_70; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_72 = 7'h42 == _GEN_793 ? L0Memory_66 : _GEN_71; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_73 = 7'h43 == _GEN_793 ? L0Memory_67 : _GEN_72; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_74 = 7'h44 == _GEN_793 ? L0Memory_68 : _GEN_73; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_75 = 7'h45 == _GEN_793 ? L0Memory_69 : _GEN_74; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_76 = 7'h46 == _GEN_793 ? L0Memory_70 : _GEN_75; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_77 = 7'h47 == _GEN_793 ? L0Memory_71 : _GEN_76; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_78 = 7'h48 == _GEN_793 ? L0Memory_72 : _GEN_77; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_79 = 7'h49 == _GEN_793 ? L0Memory_73 : _GEN_78; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_80 = 7'h4a == _GEN_793 ? L0Memory_74 : _GEN_79; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_81 = 7'h4b == _GEN_793 ? L0Memory_75 : _GEN_80; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_82 = 7'h4c == _GEN_793 ? L0Memory_76 : _GEN_81; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_83 = 7'h4d == _GEN_793 ? L0Memory_77 : _GEN_82; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_84 = 7'h4e == _GEN_793 ? L0Memory_78 : _GEN_83; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_85 = 7'h4f == _GEN_793 ? L0Memory_79 : _GEN_84; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_86 = 7'h50 == _GEN_793 ? L0Memory_80 : _GEN_85; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_87 = 7'h51 == _GEN_793 ? L0Memory_81 : _GEN_86; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_88 = 7'h52 == _GEN_793 ? L0Memory_82 : _GEN_87; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_89 = 7'h53 == _GEN_793 ? L0Memory_83 : _GEN_88; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_90 = 7'h54 == _GEN_793 ? L0Memory_84 : _GEN_89; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_91 = 7'h55 == _GEN_793 ? L0Memory_85 : _GEN_90; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_92 = 7'h56 == _GEN_793 ? L0Memory_86 : _GEN_91; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_93 = 7'h57 == _GEN_793 ? L0Memory_87 : _GEN_92; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_94 = 7'h58 == _GEN_793 ? L0Memory_88 : _GEN_93; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_95 = 7'h59 == _GEN_793 ? L0Memory_89 : _GEN_94; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_96 = 7'h5a == _GEN_793 ? L0Memory_90 : _GEN_95; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_97 = 7'h5b == _GEN_793 ? L0Memory_91 : _GEN_96; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_98 = 7'h5c == _GEN_793 ? L0Memory_92 : _GEN_97; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_99 = 7'h5d == _GEN_793 ? L0Memory_93 : _GEN_98; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_100 = 7'h5e == _GEN_793 ? L0Memory_94 : _GEN_99; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_101 = 7'h5f == _GEN_793 ? L0Memory_95 : _GEN_100; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_102 = 7'h60 == _GEN_793 ? L0Memory_96 : _GEN_101; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_103 = 7'h61 == _GEN_793 ? L0Memory_97 : _GEN_102; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_104 = 7'h62 == _GEN_793 ? L0Memory_98 : _GEN_103; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_105 = 7'h63 == _GEN_793 ? L0Memory_99 : _GEN_104; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire  _GEN_575 = _T_12 ? 1'h0 : _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 157:12]
  wire  sel5 = _T_3 ? 1'h0 : _GEN_575; // @[Conditional.scala 40:58 PEArray.scala 112:12]
  reg [15:0] mux2out_reg; // @[PEArray.scala 90:28]
  reg [15:0] mux3out_reg; // @[PEArray.scala 91:28]
  reg [9:0] count; // @[PEArray.scala 101:22]
  reg [5:0] GRU_out_width; // @[PEArray.scala 104:26]
  wire [7:0] _GEN_118 = io_control_signal_mask[8] ? 8'h0 : {{2'd0}, GRU_out_width}; // @[PEArray.scala 116:57 PEArray.scala 145:23 PEArray.scala 104:26]
  wire [9:0] _count_T_1 = count + 10'h1; // @[PEArray.scala 162:24]
  wire [9:0] _GEN_120 = count != 10'h33 ? _count_T_1 : count; // @[PEArray.scala 161:27 PEArray.scala 162:15 PEArray.scala 101:22]
  wire [9:0] _GEN_124 = count != 10'h188 ? _count_T_1 : count; // @[PEArray.scala 183:28 PEArray.scala 184:15 PEArray.scala 101:22]
  wire [9:0] _GEN_125 = count == 10'h188 ? 10'h0 : _GEN_124; // @[PEArray.scala 186:28 PEArray.scala 187:15]
  wire [2:0] _GEN_126 = count == 10'h188 ? 3'h0 : state; // @[PEArray.scala 186:28 PEArray.scala 188:15 PEArray.scala 100:22]
  wire [9:0] _GEN_127 = count != 10'h0 ? _count_T_1 : count; // @[PEArray.scala 192:32 PEArray.scala 193:15 PEArray.scala 101:22]
  wire  _T_24 = count == 10'h0; // @[PEArray.scala 195:18]
  wire [5:0] _GEN_128 = count == 10'h0 ? 6'h0 : L0Index; // @[PEArray.scala 195:26 PEArray.scala 196:17 PEArray.scala 39:24]
  wire [9:0] _T_27 = 10'h0 - 10'h1; // @[PEArray.scala 198:51]
  wire [15:0] _GEN_129 = 6'h0 == L0Index ? io_FromL1 : L0Memory_0; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_130 = 6'h1 == L0Index ? io_FromL1 : L0Memory_1; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_131 = 6'h2 == L0Index ? io_FromL1 : L0Memory_2; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_132 = 6'h3 == L0Index ? io_FromL1 : L0Memory_3; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_133 = 6'h4 == L0Index ? io_FromL1 : L0Memory_4; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_134 = 6'h5 == L0Index ? io_FromL1 : L0Memory_5; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_135 = 6'h6 == L0Index ? io_FromL1 : L0Memory_6; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_136 = 6'h7 == L0Index ? io_FromL1 : L0Memory_7; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_137 = 6'h8 == L0Index ? io_FromL1 : L0Memory_8; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_138 = 6'h9 == L0Index ? io_FromL1 : L0Memory_9; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_139 = 6'ha == L0Index ? io_FromL1 : L0Memory_10; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_140 = 6'hb == L0Index ? io_FromL1 : L0Memory_11; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_141 = 6'hc == L0Index ? io_FromL1 : L0Memory_12; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_142 = 6'hd == L0Index ? io_FromL1 : L0Memory_13; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_143 = 6'he == L0Index ? io_FromL1 : L0Memory_14; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_144 = 6'hf == L0Index ? io_FromL1 : L0Memory_15; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_145 = 6'h10 == L0Index ? io_FromL1 : L0Memory_16; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_146 = 6'h11 == L0Index ? io_FromL1 : L0Memory_17; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_147 = 6'h12 == L0Index ? io_FromL1 : L0Memory_18; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_148 = 6'h13 == L0Index ? io_FromL1 : L0Memory_19; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_149 = 6'h14 == L0Index ? io_FromL1 : L0Memory_20; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_150 = 6'h15 == L0Index ? io_FromL1 : L0Memory_21; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_151 = 6'h16 == L0Index ? io_FromL1 : L0Memory_22; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_152 = 6'h17 == L0Index ? io_FromL1 : L0Memory_23; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_153 = 6'h18 == L0Index ? io_FromL1 : L0Memory_24; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_154 = 6'h19 == L0Index ? io_FromL1 : L0Memory_25; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_155 = 6'h1a == L0Index ? io_FromL1 : L0Memory_26; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_156 = 6'h1b == L0Index ? io_FromL1 : L0Memory_27; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_157 = 6'h1c == L0Index ? io_FromL1 : L0Memory_28; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_158 = 6'h1d == L0Index ? io_FromL1 : L0Memory_29; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_159 = 6'h1e == L0Index ? io_FromL1 : L0Memory_30; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_160 = 6'h1f == L0Index ? io_FromL1 : L0Memory_31; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_161 = 6'h20 == L0Index ? io_FromL1 : L0Memory_32; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_162 = 6'h21 == L0Index ? io_FromL1 : L0Memory_33; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_163 = 6'h22 == L0Index ? io_FromL1 : L0Memory_34; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_164 = 6'h23 == L0Index ? io_FromL1 : L0Memory_35; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_165 = 6'h24 == L0Index ? io_FromL1 : L0Memory_36; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_166 = 6'h25 == L0Index ? io_FromL1 : L0Memory_37; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_167 = 6'h26 == L0Index ? io_FromL1 : L0Memory_38; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_168 = 6'h27 == L0Index ? io_FromL1 : L0Memory_39; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_169 = 6'h28 == L0Index ? io_FromL1 : L0Memory_40; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_170 = 6'h29 == L0Index ? io_FromL1 : L0Memory_41; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_171 = 6'h2a == L0Index ? io_FromL1 : L0Memory_42; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_172 = 6'h2b == L0Index ? io_FromL1 : L0Memory_43; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_173 = 6'h2c == L0Index ? io_FromL1 : L0Memory_44; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_174 = 6'h2d == L0Index ? io_FromL1 : L0Memory_45; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_175 = 6'h2e == L0Index ? io_FromL1 : L0Memory_46; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_176 = 6'h2f == L0Index ? io_FromL1 : L0Memory_47; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_177 = 6'h30 == L0Index ? io_FromL1 : L0Memory_48; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_178 = 6'h31 == L0Index ? io_FromL1 : L0Memory_49; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_179 = 6'h32 == L0Index ? io_FromL1 : L0Memory_50; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_180 = 6'h33 == L0Index ? io_FromL1 : L0Memory_51; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_181 = 6'h34 == L0Index ? io_FromL1 : L0Memory_52; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_182 = 6'h35 == L0Index ? io_FromL1 : L0Memory_53; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_183 = 6'h36 == L0Index ? io_FromL1 : L0Memory_54; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_184 = 6'h37 == L0Index ? io_FromL1 : L0Memory_55; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_185 = 6'h38 == L0Index ? io_FromL1 : L0Memory_56; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_186 = 6'h39 == L0Index ? io_FromL1 : L0Memory_57; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_187 = 6'h3a == L0Index ? io_FromL1 : L0Memory_58; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_188 = 6'h3b == L0Index ? io_FromL1 : L0Memory_59; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_189 = 6'h3c == L0Index ? io_FromL1 : L0Memory_60; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_190 = 6'h3d == L0Index ? io_FromL1 : L0Memory_61; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_191 = 6'h3e == L0Index ? io_FromL1 : L0Memory_62; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_192 = 6'h3f == L0Index ? io_FromL1 : L0Memory_63; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_193 = 7'h40 == _GEN_793 ? io_FromL1 : L0Memory_64; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_194 = 7'h41 == _GEN_793 ? io_FromL1 : L0Memory_65; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_195 = 7'h42 == _GEN_793 ? io_FromL1 : L0Memory_66; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_196 = 7'h43 == _GEN_793 ? io_FromL1 : L0Memory_67; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_197 = 7'h44 == _GEN_793 ? io_FromL1 : L0Memory_68; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_198 = 7'h45 == _GEN_793 ? io_FromL1 : L0Memory_69; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_199 = 7'h46 == _GEN_793 ? io_FromL1 : L0Memory_70; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_200 = 7'h47 == _GEN_793 ? io_FromL1 : L0Memory_71; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_201 = 7'h48 == _GEN_793 ? io_FromL1 : L0Memory_72; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_202 = 7'h49 == _GEN_793 ? io_FromL1 : L0Memory_73; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_203 = 7'h4a == _GEN_793 ? io_FromL1 : L0Memory_74; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_204 = 7'h4b == _GEN_793 ? io_FromL1 : L0Memory_75; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_205 = 7'h4c == _GEN_793 ? io_FromL1 : L0Memory_76; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_206 = 7'h4d == _GEN_793 ? io_FromL1 : L0Memory_77; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_207 = 7'h4e == _GEN_793 ? io_FromL1 : L0Memory_78; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_208 = 7'h4f == _GEN_793 ? io_FromL1 : L0Memory_79; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_209 = 7'h50 == _GEN_793 ? io_FromL1 : L0Memory_80; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_210 = 7'h51 == _GEN_793 ? io_FromL1 : L0Memory_81; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_211 = 7'h52 == _GEN_793 ? io_FromL1 : L0Memory_82; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_212 = 7'h53 == _GEN_793 ? io_FromL1 : L0Memory_83; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_213 = 7'h54 == _GEN_793 ? io_FromL1 : L0Memory_84; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_214 = 7'h55 == _GEN_793 ? io_FromL1 : L0Memory_85; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_215 = 7'h56 == _GEN_793 ? io_FromL1 : L0Memory_86; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_216 = 7'h57 == _GEN_793 ? io_FromL1 : L0Memory_87; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_217 = 7'h58 == _GEN_793 ? io_FromL1 : L0Memory_88; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_218 = 7'h59 == _GEN_793 ? io_FromL1 : L0Memory_89; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_219 = 7'h5a == _GEN_793 ? io_FromL1 : L0Memory_90; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_220 = 7'h5b == _GEN_793 ? io_FromL1 : L0Memory_91; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_221 = 7'h5c == _GEN_793 ? io_FromL1 : L0Memory_92; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_222 = 7'h5d == _GEN_793 ? io_FromL1 : L0Memory_93; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_223 = 7'h5e == _GEN_793 ? io_FromL1 : L0Memory_94; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_224 = 7'h5f == _GEN_793 ? io_FromL1 : L0Memory_95; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_225 = 7'h60 == _GEN_793 ? io_FromL1 : L0Memory_96; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_226 = 7'h61 == _GEN_793 ? io_FromL1 : L0Memory_97; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_227 = 7'h62 == _GEN_793 ? io_FromL1 : L0Memory_98; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_228 = 7'h63 == _GEN_793 ? io_FromL1 : L0Memory_99; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [5:0] _L0Index_T_2 = L0Index + 6'h1; // @[PEArray.scala 200:28]
  wire [15:0] _GEN_229 = count >= 10'h1 & count <= _T_27 ? _GEN_129 : L0Memory_0; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_230 = count >= 10'h1 & count <= _T_27 ? _GEN_130 : L0Memory_1; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_231 = count >= 10'h1 & count <= _T_27 ? _GEN_131 : L0Memory_2; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_232 = count >= 10'h1 & count <= _T_27 ? _GEN_132 : L0Memory_3; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_233 = count >= 10'h1 & count <= _T_27 ? _GEN_133 : L0Memory_4; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_234 = count >= 10'h1 & count <= _T_27 ? _GEN_134 : L0Memory_5; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_235 = count >= 10'h1 & count <= _T_27 ? _GEN_135 : L0Memory_6; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_236 = count >= 10'h1 & count <= _T_27 ? _GEN_136 : L0Memory_7; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_237 = count >= 10'h1 & count <= _T_27 ? _GEN_137 : L0Memory_8; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_238 = count >= 10'h1 & count <= _T_27 ? _GEN_138 : L0Memory_9; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_239 = count >= 10'h1 & count <= _T_27 ? _GEN_139 : L0Memory_10; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_240 = count >= 10'h1 & count <= _T_27 ? _GEN_140 : L0Memory_11; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_241 = count >= 10'h1 & count <= _T_27 ? _GEN_141 : L0Memory_12; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_242 = count >= 10'h1 & count <= _T_27 ? _GEN_142 : L0Memory_13; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_243 = count >= 10'h1 & count <= _T_27 ? _GEN_143 : L0Memory_14; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_244 = count >= 10'h1 & count <= _T_27 ? _GEN_144 : L0Memory_15; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_245 = count >= 10'h1 & count <= _T_27 ? _GEN_145 : L0Memory_16; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_246 = count >= 10'h1 & count <= _T_27 ? _GEN_146 : L0Memory_17; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_247 = count >= 10'h1 & count <= _T_27 ? _GEN_147 : L0Memory_18; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_248 = count >= 10'h1 & count <= _T_27 ? _GEN_148 : L0Memory_19; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_249 = count >= 10'h1 & count <= _T_27 ? _GEN_149 : L0Memory_20; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_250 = count >= 10'h1 & count <= _T_27 ? _GEN_150 : L0Memory_21; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_251 = count >= 10'h1 & count <= _T_27 ? _GEN_151 : L0Memory_22; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_252 = count >= 10'h1 & count <= _T_27 ? _GEN_152 : L0Memory_23; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_253 = count >= 10'h1 & count <= _T_27 ? _GEN_153 : L0Memory_24; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_254 = count >= 10'h1 & count <= _T_27 ? _GEN_154 : L0Memory_25; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_255 = count >= 10'h1 & count <= _T_27 ? _GEN_155 : L0Memory_26; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_256 = count >= 10'h1 & count <= _T_27 ? _GEN_156 : L0Memory_27; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_257 = count >= 10'h1 & count <= _T_27 ? _GEN_157 : L0Memory_28; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_258 = count >= 10'h1 & count <= _T_27 ? _GEN_158 : L0Memory_29; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_259 = count >= 10'h1 & count <= _T_27 ? _GEN_159 : L0Memory_30; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_260 = count >= 10'h1 & count <= _T_27 ? _GEN_160 : L0Memory_31; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_261 = count >= 10'h1 & count <= _T_27 ? _GEN_161 : L0Memory_32; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_262 = count >= 10'h1 & count <= _T_27 ? _GEN_162 : L0Memory_33; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_263 = count >= 10'h1 & count <= _T_27 ? _GEN_163 : L0Memory_34; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_264 = count >= 10'h1 & count <= _T_27 ? _GEN_164 : L0Memory_35; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_265 = count >= 10'h1 & count <= _T_27 ? _GEN_165 : L0Memory_36; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_266 = count >= 10'h1 & count <= _T_27 ? _GEN_166 : L0Memory_37; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_267 = count >= 10'h1 & count <= _T_27 ? _GEN_167 : L0Memory_38; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_268 = count >= 10'h1 & count <= _T_27 ? _GEN_168 : L0Memory_39; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_269 = count >= 10'h1 & count <= _T_27 ? _GEN_169 : L0Memory_40; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_270 = count >= 10'h1 & count <= _T_27 ? _GEN_170 : L0Memory_41; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_271 = count >= 10'h1 & count <= _T_27 ? _GEN_171 : L0Memory_42; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_272 = count >= 10'h1 & count <= _T_27 ? _GEN_172 : L0Memory_43; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_273 = count >= 10'h1 & count <= _T_27 ? _GEN_173 : L0Memory_44; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_274 = count >= 10'h1 & count <= _T_27 ? _GEN_174 : L0Memory_45; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_275 = count >= 10'h1 & count <= _T_27 ? _GEN_175 : L0Memory_46; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_276 = count >= 10'h1 & count <= _T_27 ? _GEN_176 : L0Memory_47; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_277 = count >= 10'h1 & count <= _T_27 ? _GEN_177 : L0Memory_48; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_278 = count >= 10'h1 & count <= _T_27 ? _GEN_178 : L0Memory_49; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_279 = count >= 10'h1 & count <= _T_27 ? _GEN_179 : L0Memory_50; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_280 = count >= 10'h1 & count <= _T_27 ? _GEN_180 : L0Memory_51; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_281 = count >= 10'h1 & count <= _T_27 ? _GEN_181 : L0Memory_52; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_282 = count >= 10'h1 & count <= _T_27 ? _GEN_182 : L0Memory_53; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_283 = count >= 10'h1 & count <= _T_27 ? _GEN_183 : L0Memory_54; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_284 = count >= 10'h1 & count <= _T_27 ? _GEN_184 : L0Memory_55; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_285 = count >= 10'h1 & count <= _T_27 ? _GEN_185 : L0Memory_56; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_286 = count >= 10'h1 & count <= _T_27 ? _GEN_186 : L0Memory_57; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_287 = count >= 10'h1 & count <= _T_27 ? _GEN_187 : L0Memory_58; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_288 = count >= 10'h1 & count <= _T_27 ? _GEN_188 : L0Memory_59; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_289 = count >= 10'h1 & count <= _T_27 ? _GEN_189 : L0Memory_60; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_290 = count >= 10'h1 & count <= _T_27 ? _GEN_190 : L0Memory_61; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_291 = count >= 10'h1 & count <= _T_27 ? _GEN_191 : L0Memory_62; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_292 = count >= 10'h1 & count <= _T_27 ? _GEN_192 : L0Memory_63; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_293 = count >= 10'h1 & count <= _T_27 ? _GEN_193 : L0Memory_64; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_294 = count >= 10'h1 & count <= _T_27 ? _GEN_194 : L0Memory_65; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_295 = count >= 10'h1 & count <= _T_27 ? _GEN_195 : L0Memory_66; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_296 = count >= 10'h1 & count <= _T_27 ? _GEN_196 : L0Memory_67; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_297 = count >= 10'h1 & count <= _T_27 ? _GEN_197 : L0Memory_68; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_298 = count >= 10'h1 & count <= _T_27 ? _GEN_198 : L0Memory_69; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_299 = count >= 10'h1 & count <= _T_27 ? _GEN_199 : L0Memory_70; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_300 = count >= 10'h1 & count <= _T_27 ? _GEN_200 : L0Memory_71; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_301 = count >= 10'h1 & count <= _T_27 ? _GEN_201 : L0Memory_72; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_302 = count >= 10'h1 & count <= _T_27 ? _GEN_202 : L0Memory_73; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_303 = count >= 10'h1 & count <= _T_27 ? _GEN_203 : L0Memory_74; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_304 = count >= 10'h1 & count <= _T_27 ? _GEN_204 : L0Memory_75; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_305 = count >= 10'h1 & count <= _T_27 ? _GEN_205 : L0Memory_76; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_306 = count >= 10'h1 & count <= _T_27 ? _GEN_206 : L0Memory_77; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_307 = count >= 10'h1 & count <= _T_27 ? _GEN_207 : L0Memory_78; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_308 = count >= 10'h1 & count <= _T_27 ? _GEN_208 : L0Memory_79; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_309 = count >= 10'h1 & count <= _T_27 ? _GEN_209 : L0Memory_80; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_310 = count >= 10'h1 & count <= _T_27 ? _GEN_210 : L0Memory_81; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_311 = count >= 10'h1 & count <= _T_27 ? _GEN_211 : L0Memory_82; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_312 = count >= 10'h1 & count <= _T_27 ? _GEN_212 : L0Memory_83; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_313 = count >= 10'h1 & count <= _T_27 ? _GEN_213 : L0Memory_84; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_314 = count >= 10'h1 & count <= _T_27 ? _GEN_214 : L0Memory_85; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_315 = count >= 10'h1 & count <= _T_27 ? _GEN_215 : L0Memory_86; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_316 = count >= 10'h1 & count <= _T_27 ? _GEN_216 : L0Memory_87; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_317 = count >= 10'h1 & count <= _T_27 ? _GEN_217 : L0Memory_88; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_318 = count >= 10'h1 & count <= _T_27 ? _GEN_218 : L0Memory_89; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_319 = count >= 10'h1 & count <= _T_27 ? _GEN_219 : L0Memory_90; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_320 = count >= 10'h1 & count <= _T_27 ? _GEN_220 : L0Memory_91; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_321 = count >= 10'h1 & count <= _T_27 ? _GEN_221 : L0Memory_92; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_322 = count >= 10'h1 & count <= _T_27 ? _GEN_222 : L0Memory_93; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_323 = count >= 10'h1 & count <= _T_27 ? _GEN_223 : L0Memory_94; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_324 = count >= 10'h1 & count <= _T_27 ? _GEN_224 : L0Memory_95; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_325 = count >= 10'h1 & count <= _T_27 ? _GEN_225 : L0Memory_96; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_326 = count >= 10'h1 & count <= _T_27 ? _GEN_226 : L0Memory_97; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_327 = count >= 10'h1 & count <= _T_27 ? _GEN_227 : L0Memory_98; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_328 = count >= 10'h1 & count <= _T_27 ? _GEN_228 : L0Memory_99; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [5:0] _GEN_329 = count >= 10'h1 & count <= _T_27 ? _L0Index_T_2 : _GEN_128; // @[PEArray.scala 198:59 PEArray.scala 200:17]
  wire [9:0] _GEN_330 = _T_24 ? 10'h0 : _GEN_127; // @[PEArray.scala 202:32 PEArray.scala 203:15]
  wire [2:0] _GEN_331 = _T_24 ? 3'h0 : state; // @[PEArray.scala 202:32 PEArray.scala 204:15 PEArray.scala 100:22]
  wire [9:0] _GEN_865 = {{4'd0}, GRU_out_width}; // @[PEArray.scala 220:19]
  wire [9:0] _GEN_0 = count % _GEN_865; // @[PEArray.scala 220:19]
  wire [5:0] _T_36 = _GEN_0[5:0]; // @[PEArray.scala 220:19]
  wire [5:0] _T_38 = GRU_out_width - 6'h1; // @[PEArray.scala 220:55]
  wire [5:0] _GEN_334 = _T_36 == _T_38 ? _L0Index_T_2 : 6'h0; // @[PEArray.scala 220:62 PEArray.scala 221:17 PEArray.scala 214:15]
  wire [5:0] _GEN_346 = _T_41 ? _GEN_334 : L0Index; // @[Conditional.scala 39:67 PEArray.scala 39:24]
  wire [9:0] _GEN_347 = _T_41 ? _GEN_330 : count; // @[Conditional.scala 39:67 PEArray.scala 101:22]
  wire [2:0] _GEN_348 = _T_41 ? _GEN_331 : state; // @[Conditional.scala 39:67 PEArray.scala 100:22]
  wire [5:0] _GEN_353 = _T_31 ? _GEN_334 : _GEN_346; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_354 = _T_31 ? _GEN_330 : _GEN_347; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_355 = _T_31 ? _GEN_331 : _GEN_348; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_356 = _T_22 ? _GEN_330 : _GEN_354; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_357 = _T_22 ? _GEN_329 : _GEN_353; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_458 = _T_22 ? _GEN_331 : _GEN_355; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_690 = _T_3 ? _GEN_118 : {{2'd0}, GRU_out_width}; // @[Conditional.scala 40:58 PEArray.scala 104:26]
  FP16MulAdder FP16MAC ( // @[PEArray.scala 72:23]
    .io_a(FP16MAC_io_a),
    .io_b(FP16MAC_io_b),
    .io_c(FP16MAC_io_c),
    .io_out(FP16MAC_io_out)
  );
  assign io_ToRightPE = mux3out_reg; // @[PEArray.scala 95:16]
  assign io_ToBelowPE = mux2out_reg; // @[PEArray.scala 94:16]
  assign FP16MAC_io_a = sel1 ? io_FromL1 : io_FromLeftPE; // @[PEArray.scala 50:14 PEArray.scala 50:23 PEArray.scala 51:24]
  assign FP16MAC_io_b = sel5 ? mux4out : _GEN_105; // @[PEArray.scala 77:13 PEArray.scala 78:18 PEArray.scala 81:18]
  assign FP16MAC_io_c = sel5 ? _GEN_105 : mux4out; // @[PEArray.scala 77:13 PEArray.scala 79:18 PEArray.scala 82:18]
  always @(posedge clock) begin
    if (reset) begin // @[PEArray.scala 39:24]
      L0Index <= 6'h0; // @[PEArray.scala 39:24]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h0; // @[PEArray.scala 159:15]
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h6; // @[PEArray.scala 181:15]
      end else begin
        L0Index <= _GEN_357;
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_0 <= _GEN_229;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_1 <= _GEN_230;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_2 <= _GEN_231;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_3 <= _GEN_232;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_4 <= _GEN_233;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_5 <= _GEN_234;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_6 <= _GEN_235;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_7 <= _GEN_236;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_8 <= _GEN_237;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_9 <= _GEN_238;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_10 <= _GEN_239;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_11 <= _GEN_240;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_12 <= _GEN_241;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_13 <= _GEN_242;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_14 <= _GEN_243;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_15 <= _GEN_244;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_16 <= _GEN_245;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_17 <= _GEN_246;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_18 <= _GEN_247;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_19 <= _GEN_248;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_20 <= _GEN_249;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_21 <= _GEN_250;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_22 <= _GEN_251;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_23 <= _GEN_252;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_24 <= _GEN_253;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_25 <= _GEN_254;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_26 <= _GEN_255;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_27 <= _GEN_256;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_28 <= _GEN_257;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_29 <= _GEN_258;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_30 <= _GEN_259;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_31 <= _GEN_260;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_32 <= _GEN_261;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_33 <= _GEN_262;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_34 <= _GEN_263;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_35 <= _GEN_264;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_36 <= _GEN_265;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_37 <= _GEN_266;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_38 <= _GEN_267;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_39 <= _GEN_268;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_40 <= _GEN_269;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_41 <= _GEN_270;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_42 <= _GEN_271;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_43 <= _GEN_272;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_44 <= _GEN_273;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_45 <= _GEN_274;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_46 <= _GEN_275;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_47 <= _GEN_276;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_48 <= _GEN_277;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_49 <= _GEN_278;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_50 <= _GEN_279;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_51 <= _GEN_280;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_52 <= _GEN_281;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_53 <= _GEN_282;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_54 <= _GEN_283;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_55 <= _GEN_284;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_56 <= _GEN_285;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_57 <= _GEN_286;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_58 <= _GEN_287;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_59 <= _GEN_288;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_60 <= _GEN_289;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_61 <= _GEN_290;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_62 <= _GEN_291;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_63 <= _GEN_292;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_64 <= _GEN_293;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_65 <= _GEN_294;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_66 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_67 <= _GEN_296;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_68 <= _GEN_297;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_69 <= _GEN_298;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_70 <= _GEN_299;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_71 <= _GEN_300;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_72 <= _GEN_301;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_73 <= _GEN_302;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_74 <= _GEN_303;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_75 <= _GEN_304;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_76 <= _GEN_305;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_77 <= _GEN_306;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_78 <= _GEN_307;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_79 <= _GEN_308;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_80 <= _GEN_309;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_81 <= _GEN_310;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_82 <= _GEN_311;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_83 <= _GEN_312;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_84 <= _GEN_313;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_85 <= _GEN_314;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_86 <= _GEN_315;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_87 <= _GEN_316;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_88 <= _GEN_317;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_89 <= _GEN_318;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_90 <= _GEN_319;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_91 <= _GEN_320;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_92 <= _GEN_321;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_93 <= _GEN_322;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_94 <= _GEN_323;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_95 <= _GEN_324;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_96 <= _GEN_325;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_97 <= _GEN_326;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_98 <= _GEN_327;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_99 <= _GEN_328;
          end
        end
      end
    end
    if (reset) begin // @[PEArray.scala 100:22]
      state <= 3'h0; // @[PEArray.scala 100:22]
    end else if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[8]) begin // @[PEArray.scala 116:57]
        state <= 3'h1;
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      if (count == 10'h33) begin // @[PEArray.scala 164:27]
        state <= 3'h0; // @[PEArray.scala 166:15]
      end
    end else if (_T_16) begin // @[Conditional.scala 39:67]
      state <= _GEN_126;
    end else begin
      state <= _GEN_458;
    end
    if (reset) begin // @[PEArray.scala 90:28]
      mux2out_reg <= 16'h0; // @[PEArray.scala 90:28]
    end else begin
      mux2out_reg <= MAC_out; // @[PEArray.scala 90:28]
    end
    if (reset) begin // @[PEArray.scala 91:28]
      mux3out_reg <= 16'h0; // @[PEArray.scala 91:28]
    end else if (sel3) begin // @[PEArray.scala 56:14]
      mux3out_reg <= MAC_out; // @[PEArray.scala 56:23]
    end else if (sel1) begin // @[PEArray.scala 50:14]
      mux3out_reg <= io_FromL1; // @[PEArray.scala 50:23]
    end else begin
      mux3out_reg <= io_FromLeftPE; // @[PEArray.scala 51:24]
    end
    if (reset) begin // @[PEArray.scala 101:22]
      count <= 10'h0; // @[PEArray.scala 101:22]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        if (count == 10'h33) begin // @[PEArray.scala 164:27]
          count <= 10'h0; // @[PEArray.scala 165:15]
        end else begin
          count <= _GEN_120;
        end
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        count <= _GEN_125;
      end else begin
        count <= _GEN_356;
      end
    end
    GRU_out_width <= _GEN_690[5:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  L0Index = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  L0Memory_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  L0Memory_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  L0Memory_2 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  L0Memory_3 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  L0Memory_4 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  L0Memory_5 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  L0Memory_6 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  L0Memory_7 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  L0Memory_8 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  L0Memory_9 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  L0Memory_10 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  L0Memory_11 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  L0Memory_12 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  L0Memory_13 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  L0Memory_14 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  L0Memory_15 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  L0Memory_16 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  L0Memory_17 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  L0Memory_18 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  L0Memory_19 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  L0Memory_20 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  L0Memory_21 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  L0Memory_22 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  L0Memory_23 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  L0Memory_24 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  L0Memory_25 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  L0Memory_26 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  L0Memory_27 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  L0Memory_28 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  L0Memory_29 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  L0Memory_30 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  L0Memory_31 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  L0Memory_32 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  L0Memory_33 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  L0Memory_34 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  L0Memory_35 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  L0Memory_36 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  L0Memory_37 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  L0Memory_38 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  L0Memory_39 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  L0Memory_40 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  L0Memory_41 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  L0Memory_42 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  L0Memory_43 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  L0Memory_44 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  L0Memory_45 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  L0Memory_46 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  L0Memory_47 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  L0Memory_48 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  L0Memory_49 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  L0Memory_50 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  L0Memory_51 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  L0Memory_52 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  L0Memory_53 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  L0Memory_54 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  L0Memory_55 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  L0Memory_56 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  L0Memory_57 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  L0Memory_58 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  L0Memory_59 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  L0Memory_60 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  L0Memory_61 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  L0Memory_62 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  L0Memory_63 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  L0Memory_64 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  L0Memory_65 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  L0Memory_66 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  L0Memory_67 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  L0Memory_68 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  L0Memory_69 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  L0Memory_70 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  L0Memory_71 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  L0Memory_72 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  L0Memory_73 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  L0Memory_74 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  L0Memory_75 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  L0Memory_76 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  L0Memory_77 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  L0Memory_78 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  L0Memory_79 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  L0Memory_80 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  L0Memory_81 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  L0Memory_82 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  L0Memory_83 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  L0Memory_84 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  L0Memory_85 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  L0Memory_86 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  L0Memory_87 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  L0Memory_88 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  L0Memory_89 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  L0Memory_90 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  L0Memory_91 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  L0Memory_92 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  L0Memory_93 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  L0Memory_94 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  L0Memory_95 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  L0Memory_96 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  L0Memory_97 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  L0Memory_98 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  L0Memory_99 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  state = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  mux2out_reg = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  mux3out_reg = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  count = _RAND_104[9:0];
  _RAND_105 = {1{`RANDOM}};
  GRU_out_width = _RAND_105[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PE_10(
  input         clock,
  input         reset,
  input  [15:0] io_FromAbovePE,
  input  [15:0] io_FromLeftPE,
  input  [15:0] io_FromL1,
  input  [11:0] io_control_signal_mask,
  output [15:0] io_ToRightPE,
  output [15:0] io_ToBelowPE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] FP16MAC_io_a; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_b; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_c; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_out; // @[PEArray.scala 72:23]
  reg [5:0] L0Index; // @[PEArray.scala 39:24]
  reg [15:0] L0Memory_0; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_1; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_2; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_3; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_4; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_5; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_6; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_7; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_8; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_9; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_10; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_11; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_12; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_13; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_14; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_15; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_16; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_17; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_18; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_19; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_20; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_21; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_22; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_23; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_24; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_25; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_26; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_27; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_28; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_29; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_30; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_31; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_32; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_33; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_34; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_35; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_36; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_37; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_38; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_39; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_40; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_41; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_42; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_43; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_44; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_45; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_46; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_47; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_48; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_49; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_50; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_51; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_52; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_53; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_54; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_55; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_56; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_57; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_58; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_59; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_60; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_61; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_62; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_63; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_64; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_65; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_66; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_67; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_68; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_69; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_70; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_71; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_72; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_73; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_74; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_75; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_76; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_77; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_78; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_79; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_80; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_81; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_82; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_83; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_84; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_85; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_86; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_87; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_88; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_89; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_90; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_91; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_92; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_93; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_94; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_95; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_96; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_97; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_98; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_99; // @[PEArray.scala 40:21]
  reg [2:0] state; // @[PEArray.scala 100:22]
  wire  _T_3 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_12 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_16 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_22 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_31 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_41 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_342 = _T_41 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 231:12 PEArray.scala 32:8]
  wire  _GEN_349 = _T_31 ? 1'h0 : _GEN_342; // @[Conditional.scala 39:67 PEArray.scala 208:12]
  wire  _GEN_459 = _T_22 | _GEN_349; // @[Conditional.scala 39:67 PEArray.scala 32:8]
  wire  _GEN_463 = _T_16 ? 1'h0 : _GEN_459; // @[Conditional.scala 39:67]
  wire  _GEN_572 = _T_12 | _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 149:12]
  wire  sel1 = _T_3 | _GEN_572; // @[Conditional.scala 40:58 PEArray.scala 108:12]
  wire [15:0] MAC_out = FP16MAC_io_out; // @[PEArray.scala 47:21 PEArray.scala 85:11]
  wire  _GEN_465 = _T_16 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 177:12]
  wire  _GEN_580 = _T_12 | _GEN_465; // @[Conditional.scala 39:67 PEArray.scala 34:8]
  wire  sel3 = _T_3 | _GEN_580; // @[Conditional.scala 40:58 PEArray.scala 110:12]
  wire [1:0] _GEN_344 = _T_41 ? 2'h2 : 2'h0; // @[Conditional.scala 39:67 PEArray.scala 233:12 PEArray.scala 35:8]
  wire [1:0] _GEN_351 = _T_31 ? 2'h2 : _GEN_344; // @[Conditional.scala 39:67 PEArray.scala 210:12]
  wire [1:0] _GEN_461 = _T_22 ? 2'h0 : _GEN_351; // @[Conditional.scala 39:67 PEArray.scala 35:8]
  wire [1:0] _GEN_466 = _T_16 ? 2'h0 : _GEN_461; // @[Conditional.scala 39:67 PEArray.scala 178:12]
  wire [1:0] _GEN_574 = _T_12 ? 2'h1 : _GEN_466; // @[Conditional.scala 39:67]
  wire [1:0] sel4 = _T_3 ? 2'h0 : _GEN_574; // @[Conditional.scala 40:58 PEArray.scala 111:12]
  wire [15:0] _GEN_3 = sel4 == 2'h2 ? io_FromL1 : 16'h0; // @[PEArray.scala 65:28 PEArray.scala 66:15 PEArray.scala 69:15]
  wire [15:0] _GEN_4 = sel4 == 2'h1 ? io_FromAbovePE : _GEN_3; // @[PEArray.scala 62:28 PEArray.scala 63:15]
  wire [15:0] mux4out = sel4 == 2'h0 ? 16'h0 : _GEN_4; // @[PEArray.scala 59:22 PEArray.scala 60:13]
  wire [15:0] _GEN_7 = 6'h1 == L0Index ? L0Memory_1 : L0Memory_0; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_8 = 6'h2 == L0Index ? L0Memory_2 : _GEN_7; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_9 = 6'h3 == L0Index ? L0Memory_3 : _GEN_8; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_10 = 6'h4 == L0Index ? L0Memory_4 : _GEN_9; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_11 = 6'h5 == L0Index ? L0Memory_5 : _GEN_10; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_12 = 6'h6 == L0Index ? L0Memory_6 : _GEN_11; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_13 = 6'h7 == L0Index ? L0Memory_7 : _GEN_12; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_14 = 6'h8 == L0Index ? L0Memory_8 : _GEN_13; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_15 = 6'h9 == L0Index ? L0Memory_9 : _GEN_14; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_16 = 6'ha == L0Index ? L0Memory_10 : _GEN_15; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_17 = 6'hb == L0Index ? L0Memory_11 : _GEN_16; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_18 = 6'hc == L0Index ? L0Memory_12 : _GEN_17; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_19 = 6'hd == L0Index ? L0Memory_13 : _GEN_18; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_20 = 6'he == L0Index ? L0Memory_14 : _GEN_19; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_21 = 6'hf == L0Index ? L0Memory_15 : _GEN_20; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_22 = 6'h10 == L0Index ? L0Memory_16 : _GEN_21; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_23 = 6'h11 == L0Index ? L0Memory_17 : _GEN_22; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_24 = 6'h12 == L0Index ? L0Memory_18 : _GEN_23; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_25 = 6'h13 == L0Index ? L0Memory_19 : _GEN_24; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_26 = 6'h14 == L0Index ? L0Memory_20 : _GEN_25; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_27 = 6'h15 == L0Index ? L0Memory_21 : _GEN_26; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_28 = 6'h16 == L0Index ? L0Memory_22 : _GEN_27; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_29 = 6'h17 == L0Index ? L0Memory_23 : _GEN_28; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_30 = 6'h18 == L0Index ? L0Memory_24 : _GEN_29; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_31 = 6'h19 == L0Index ? L0Memory_25 : _GEN_30; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_32 = 6'h1a == L0Index ? L0Memory_26 : _GEN_31; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_33 = 6'h1b == L0Index ? L0Memory_27 : _GEN_32; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_34 = 6'h1c == L0Index ? L0Memory_28 : _GEN_33; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_35 = 6'h1d == L0Index ? L0Memory_29 : _GEN_34; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_36 = 6'h1e == L0Index ? L0Memory_30 : _GEN_35; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_37 = 6'h1f == L0Index ? L0Memory_31 : _GEN_36; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_38 = 6'h20 == L0Index ? L0Memory_32 : _GEN_37; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_39 = 6'h21 == L0Index ? L0Memory_33 : _GEN_38; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_40 = 6'h22 == L0Index ? L0Memory_34 : _GEN_39; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_41 = 6'h23 == L0Index ? L0Memory_35 : _GEN_40; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_42 = 6'h24 == L0Index ? L0Memory_36 : _GEN_41; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_43 = 6'h25 == L0Index ? L0Memory_37 : _GEN_42; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_44 = 6'h26 == L0Index ? L0Memory_38 : _GEN_43; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_45 = 6'h27 == L0Index ? L0Memory_39 : _GEN_44; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_46 = 6'h28 == L0Index ? L0Memory_40 : _GEN_45; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_47 = 6'h29 == L0Index ? L0Memory_41 : _GEN_46; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_48 = 6'h2a == L0Index ? L0Memory_42 : _GEN_47; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_49 = 6'h2b == L0Index ? L0Memory_43 : _GEN_48; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_50 = 6'h2c == L0Index ? L0Memory_44 : _GEN_49; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_51 = 6'h2d == L0Index ? L0Memory_45 : _GEN_50; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_52 = 6'h2e == L0Index ? L0Memory_46 : _GEN_51; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_53 = 6'h2f == L0Index ? L0Memory_47 : _GEN_52; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_54 = 6'h30 == L0Index ? L0Memory_48 : _GEN_53; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_55 = 6'h31 == L0Index ? L0Memory_49 : _GEN_54; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_56 = 6'h32 == L0Index ? L0Memory_50 : _GEN_55; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_57 = 6'h33 == L0Index ? L0Memory_51 : _GEN_56; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_58 = 6'h34 == L0Index ? L0Memory_52 : _GEN_57; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_59 = 6'h35 == L0Index ? L0Memory_53 : _GEN_58; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_60 = 6'h36 == L0Index ? L0Memory_54 : _GEN_59; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_61 = 6'h37 == L0Index ? L0Memory_55 : _GEN_60; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_62 = 6'h38 == L0Index ? L0Memory_56 : _GEN_61; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_63 = 6'h39 == L0Index ? L0Memory_57 : _GEN_62; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_64 = 6'h3a == L0Index ? L0Memory_58 : _GEN_63; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_65 = 6'h3b == L0Index ? L0Memory_59 : _GEN_64; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_66 = 6'h3c == L0Index ? L0Memory_60 : _GEN_65; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_67 = 6'h3d == L0Index ? L0Memory_61 : _GEN_66; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_68 = 6'h3e == L0Index ? L0Memory_62 : _GEN_67; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_69 = 6'h3f == L0Index ? L0Memory_63 : _GEN_68; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [6:0] _GEN_793 = {{1'd0}, L0Index}; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_70 = 7'h40 == _GEN_793 ? L0Memory_64 : _GEN_69; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_71 = 7'h41 == _GEN_793 ? L0Memory_65 : _GEN_70; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_72 = 7'h42 == _GEN_793 ? L0Memory_66 : _GEN_71; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_73 = 7'h43 == _GEN_793 ? L0Memory_67 : _GEN_72; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_74 = 7'h44 == _GEN_793 ? L0Memory_68 : _GEN_73; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_75 = 7'h45 == _GEN_793 ? L0Memory_69 : _GEN_74; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_76 = 7'h46 == _GEN_793 ? L0Memory_70 : _GEN_75; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_77 = 7'h47 == _GEN_793 ? L0Memory_71 : _GEN_76; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_78 = 7'h48 == _GEN_793 ? L0Memory_72 : _GEN_77; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_79 = 7'h49 == _GEN_793 ? L0Memory_73 : _GEN_78; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_80 = 7'h4a == _GEN_793 ? L0Memory_74 : _GEN_79; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_81 = 7'h4b == _GEN_793 ? L0Memory_75 : _GEN_80; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_82 = 7'h4c == _GEN_793 ? L0Memory_76 : _GEN_81; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_83 = 7'h4d == _GEN_793 ? L0Memory_77 : _GEN_82; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_84 = 7'h4e == _GEN_793 ? L0Memory_78 : _GEN_83; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_85 = 7'h4f == _GEN_793 ? L0Memory_79 : _GEN_84; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_86 = 7'h50 == _GEN_793 ? L0Memory_80 : _GEN_85; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_87 = 7'h51 == _GEN_793 ? L0Memory_81 : _GEN_86; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_88 = 7'h52 == _GEN_793 ? L0Memory_82 : _GEN_87; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_89 = 7'h53 == _GEN_793 ? L0Memory_83 : _GEN_88; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_90 = 7'h54 == _GEN_793 ? L0Memory_84 : _GEN_89; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_91 = 7'h55 == _GEN_793 ? L0Memory_85 : _GEN_90; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_92 = 7'h56 == _GEN_793 ? L0Memory_86 : _GEN_91; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_93 = 7'h57 == _GEN_793 ? L0Memory_87 : _GEN_92; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_94 = 7'h58 == _GEN_793 ? L0Memory_88 : _GEN_93; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_95 = 7'h59 == _GEN_793 ? L0Memory_89 : _GEN_94; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_96 = 7'h5a == _GEN_793 ? L0Memory_90 : _GEN_95; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_97 = 7'h5b == _GEN_793 ? L0Memory_91 : _GEN_96; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_98 = 7'h5c == _GEN_793 ? L0Memory_92 : _GEN_97; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_99 = 7'h5d == _GEN_793 ? L0Memory_93 : _GEN_98; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_100 = 7'h5e == _GEN_793 ? L0Memory_94 : _GEN_99; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_101 = 7'h5f == _GEN_793 ? L0Memory_95 : _GEN_100; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_102 = 7'h60 == _GEN_793 ? L0Memory_96 : _GEN_101; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_103 = 7'h61 == _GEN_793 ? L0Memory_97 : _GEN_102; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_104 = 7'h62 == _GEN_793 ? L0Memory_98 : _GEN_103; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_105 = 7'h63 == _GEN_793 ? L0Memory_99 : _GEN_104; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire  _GEN_575 = _T_12 ? 1'h0 : _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 157:12]
  wire  sel5 = _T_3 ? 1'h0 : _GEN_575; // @[Conditional.scala 40:58 PEArray.scala 112:12]
  reg [15:0] mux2out_reg; // @[PEArray.scala 90:28]
  reg [15:0] mux3out_reg; // @[PEArray.scala 91:28]
  reg [9:0] count; // @[PEArray.scala 101:22]
  reg [5:0] GRU_out_width; // @[PEArray.scala 104:26]
  wire [7:0] _GEN_118 = io_control_signal_mask[8] ? 8'h0 : {{2'd0}, GRU_out_width}; // @[PEArray.scala 116:57 PEArray.scala 145:23 PEArray.scala 104:26]
  wire [9:0] _count_T_1 = count + 10'h1; // @[PEArray.scala 162:24]
  wire [9:0] _GEN_120 = count != 10'h33 ? _count_T_1 : count; // @[PEArray.scala 161:27 PEArray.scala 162:15 PEArray.scala 101:22]
  wire [9:0] _GEN_124 = count != 10'h188 ? _count_T_1 : count; // @[PEArray.scala 183:28 PEArray.scala 184:15 PEArray.scala 101:22]
  wire [9:0] _GEN_125 = count == 10'h188 ? 10'h0 : _GEN_124; // @[PEArray.scala 186:28 PEArray.scala 187:15]
  wire [2:0] _GEN_126 = count == 10'h188 ? 3'h0 : state; // @[PEArray.scala 186:28 PEArray.scala 188:15 PEArray.scala 100:22]
  wire [9:0] _GEN_127 = count != 10'h0 ? _count_T_1 : count; // @[PEArray.scala 192:32 PEArray.scala 193:15 PEArray.scala 101:22]
  wire  _T_24 = count == 10'h0; // @[PEArray.scala 195:18]
  wire [5:0] _GEN_128 = count == 10'h0 ? 6'h0 : L0Index; // @[PEArray.scala 195:26 PEArray.scala 196:17 PEArray.scala 39:24]
  wire [9:0] _T_27 = 10'h0 - 10'h1; // @[PEArray.scala 198:51]
  wire [15:0] _GEN_129 = 6'h0 == L0Index ? io_FromL1 : L0Memory_0; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_130 = 6'h1 == L0Index ? io_FromL1 : L0Memory_1; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_131 = 6'h2 == L0Index ? io_FromL1 : L0Memory_2; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_132 = 6'h3 == L0Index ? io_FromL1 : L0Memory_3; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_133 = 6'h4 == L0Index ? io_FromL1 : L0Memory_4; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_134 = 6'h5 == L0Index ? io_FromL1 : L0Memory_5; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_135 = 6'h6 == L0Index ? io_FromL1 : L0Memory_6; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_136 = 6'h7 == L0Index ? io_FromL1 : L0Memory_7; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_137 = 6'h8 == L0Index ? io_FromL1 : L0Memory_8; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_138 = 6'h9 == L0Index ? io_FromL1 : L0Memory_9; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_139 = 6'ha == L0Index ? io_FromL1 : L0Memory_10; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_140 = 6'hb == L0Index ? io_FromL1 : L0Memory_11; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_141 = 6'hc == L0Index ? io_FromL1 : L0Memory_12; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_142 = 6'hd == L0Index ? io_FromL1 : L0Memory_13; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_143 = 6'he == L0Index ? io_FromL1 : L0Memory_14; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_144 = 6'hf == L0Index ? io_FromL1 : L0Memory_15; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_145 = 6'h10 == L0Index ? io_FromL1 : L0Memory_16; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_146 = 6'h11 == L0Index ? io_FromL1 : L0Memory_17; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_147 = 6'h12 == L0Index ? io_FromL1 : L0Memory_18; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_148 = 6'h13 == L0Index ? io_FromL1 : L0Memory_19; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_149 = 6'h14 == L0Index ? io_FromL1 : L0Memory_20; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_150 = 6'h15 == L0Index ? io_FromL1 : L0Memory_21; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_151 = 6'h16 == L0Index ? io_FromL1 : L0Memory_22; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_152 = 6'h17 == L0Index ? io_FromL1 : L0Memory_23; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_153 = 6'h18 == L0Index ? io_FromL1 : L0Memory_24; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_154 = 6'h19 == L0Index ? io_FromL1 : L0Memory_25; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_155 = 6'h1a == L0Index ? io_FromL1 : L0Memory_26; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_156 = 6'h1b == L0Index ? io_FromL1 : L0Memory_27; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_157 = 6'h1c == L0Index ? io_FromL1 : L0Memory_28; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_158 = 6'h1d == L0Index ? io_FromL1 : L0Memory_29; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_159 = 6'h1e == L0Index ? io_FromL1 : L0Memory_30; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_160 = 6'h1f == L0Index ? io_FromL1 : L0Memory_31; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_161 = 6'h20 == L0Index ? io_FromL1 : L0Memory_32; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_162 = 6'h21 == L0Index ? io_FromL1 : L0Memory_33; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_163 = 6'h22 == L0Index ? io_FromL1 : L0Memory_34; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_164 = 6'h23 == L0Index ? io_FromL1 : L0Memory_35; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_165 = 6'h24 == L0Index ? io_FromL1 : L0Memory_36; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_166 = 6'h25 == L0Index ? io_FromL1 : L0Memory_37; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_167 = 6'h26 == L0Index ? io_FromL1 : L0Memory_38; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_168 = 6'h27 == L0Index ? io_FromL1 : L0Memory_39; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_169 = 6'h28 == L0Index ? io_FromL1 : L0Memory_40; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_170 = 6'h29 == L0Index ? io_FromL1 : L0Memory_41; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_171 = 6'h2a == L0Index ? io_FromL1 : L0Memory_42; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_172 = 6'h2b == L0Index ? io_FromL1 : L0Memory_43; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_173 = 6'h2c == L0Index ? io_FromL1 : L0Memory_44; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_174 = 6'h2d == L0Index ? io_FromL1 : L0Memory_45; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_175 = 6'h2e == L0Index ? io_FromL1 : L0Memory_46; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_176 = 6'h2f == L0Index ? io_FromL1 : L0Memory_47; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_177 = 6'h30 == L0Index ? io_FromL1 : L0Memory_48; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_178 = 6'h31 == L0Index ? io_FromL1 : L0Memory_49; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_179 = 6'h32 == L0Index ? io_FromL1 : L0Memory_50; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_180 = 6'h33 == L0Index ? io_FromL1 : L0Memory_51; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_181 = 6'h34 == L0Index ? io_FromL1 : L0Memory_52; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_182 = 6'h35 == L0Index ? io_FromL1 : L0Memory_53; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_183 = 6'h36 == L0Index ? io_FromL1 : L0Memory_54; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_184 = 6'h37 == L0Index ? io_FromL1 : L0Memory_55; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_185 = 6'h38 == L0Index ? io_FromL1 : L0Memory_56; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_186 = 6'h39 == L0Index ? io_FromL1 : L0Memory_57; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_187 = 6'h3a == L0Index ? io_FromL1 : L0Memory_58; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_188 = 6'h3b == L0Index ? io_FromL1 : L0Memory_59; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_189 = 6'h3c == L0Index ? io_FromL1 : L0Memory_60; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_190 = 6'h3d == L0Index ? io_FromL1 : L0Memory_61; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_191 = 6'h3e == L0Index ? io_FromL1 : L0Memory_62; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_192 = 6'h3f == L0Index ? io_FromL1 : L0Memory_63; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_193 = 7'h40 == _GEN_793 ? io_FromL1 : L0Memory_64; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_194 = 7'h41 == _GEN_793 ? io_FromL1 : L0Memory_65; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_195 = 7'h42 == _GEN_793 ? io_FromL1 : L0Memory_66; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_196 = 7'h43 == _GEN_793 ? io_FromL1 : L0Memory_67; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_197 = 7'h44 == _GEN_793 ? io_FromL1 : L0Memory_68; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_198 = 7'h45 == _GEN_793 ? io_FromL1 : L0Memory_69; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_199 = 7'h46 == _GEN_793 ? io_FromL1 : L0Memory_70; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_200 = 7'h47 == _GEN_793 ? io_FromL1 : L0Memory_71; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_201 = 7'h48 == _GEN_793 ? io_FromL1 : L0Memory_72; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_202 = 7'h49 == _GEN_793 ? io_FromL1 : L0Memory_73; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_203 = 7'h4a == _GEN_793 ? io_FromL1 : L0Memory_74; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_204 = 7'h4b == _GEN_793 ? io_FromL1 : L0Memory_75; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_205 = 7'h4c == _GEN_793 ? io_FromL1 : L0Memory_76; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_206 = 7'h4d == _GEN_793 ? io_FromL1 : L0Memory_77; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_207 = 7'h4e == _GEN_793 ? io_FromL1 : L0Memory_78; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_208 = 7'h4f == _GEN_793 ? io_FromL1 : L0Memory_79; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_209 = 7'h50 == _GEN_793 ? io_FromL1 : L0Memory_80; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_210 = 7'h51 == _GEN_793 ? io_FromL1 : L0Memory_81; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_211 = 7'h52 == _GEN_793 ? io_FromL1 : L0Memory_82; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_212 = 7'h53 == _GEN_793 ? io_FromL1 : L0Memory_83; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_213 = 7'h54 == _GEN_793 ? io_FromL1 : L0Memory_84; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_214 = 7'h55 == _GEN_793 ? io_FromL1 : L0Memory_85; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_215 = 7'h56 == _GEN_793 ? io_FromL1 : L0Memory_86; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_216 = 7'h57 == _GEN_793 ? io_FromL1 : L0Memory_87; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_217 = 7'h58 == _GEN_793 ? io_FromL1 : L0Memory_88; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_218 = 7'h59 == _GEN_793 ? io_FromL1 : L0Memory_89; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_219 = 7'h5a == _GEN_793 ? io_FromL1 : L0Memory_90; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_220 = 7'h5b == _GEN_793 ? io_FromL1 : L0Memory_91; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_221 = 7'h5c == _GEN_793 ? io_FromL1 : L0Memory_92; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_222 = 7'h5d == _GEN_793 ? io_FromL1 : L0Memory_93; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_223 = 7'h5e == _GEN_793 ? io_FromL1 : L0Memory_94; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_224 = 7'h5f == _GEN_793 ? io_FromL1 : L0Memory_95; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_225 = 7'h60 == _GEN_793 ? io_FromL1 : L0Memory_96; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_226 = 7'h61 == _GEN_793 ? io_FromL1 : L0Memory_97; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_227 = 7'h62 == _GEN_793 ? io_FromL1 : L0Memory_98; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_228 = 7'h63 == _GEN_793 ? io_FromL1 : L0Memory_99; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [5:0] _L0Index_T_2 = L0Index + 6'h1; // @[PEArray.scala 200:28]
  wire [15:0] _GEN_229 = count >= 10'h1 & count <= _T_27 ? _GEN_129 : L0Memory_0; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_230 = count >= 10'h1 & count <= _T_27 ? _GEN_130 : L0Memory_1; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_231 = count >= 10'h1 & count <= _T_27 ? _GEN_131 : L0Memory_2; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_232 = count >= 10'h1 & count <= _T_27 ? _GEN_132 : L0Memory_3; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_233 = count >= 10'h1 & count <= _T_27 ? _GEN_133 : L0Memory_4; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_234 = count >= 10'h1 & count <= _T_27 ? _GEN_134 : L0Memory_5; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_235 = count >= 10'h1 & count <= _T_27 ? _GEN_135 : L0Memory_6; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_236 = count >= 10'h1 & count <= _T_27 ? _GEN_136 : L0Memory_7; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_237 = count >= 10'h1 & count <= _T_27 ? _GEN_137 : L0Memory_8; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_238 = count >= 10'h1 & count <= _T_27 ? _GEN_138 : L0Memory_9; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_239 = count >= 10'h1 & count <= _T_27 ? _GEN_139 : L0Memory_10; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_240 = count >= 10'h1 & count <= _T_27 ? _GEN_140 : L0Memory_11; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_241 = count >= 10'h1 & count <= _T_27 ? _GEN_141 : L0Memory_12; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_242 = count >= 10'h1 & count <= _T_27 ? _GEN_142 : L0Memory_13; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_243 = count >= 10'h1 & count <= _T_27 ? _GEN_143 : L0Memory_14; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_244 = count >= 10'h1 & count <= _T_27 ? _GEN_144 : L0Memory_15; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_245 = count >= 10'h1 & count <= _T_27 ? _GEN_145 : L0Memory_16; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_246 = count >= 10'h1 & count <= _T_27 ? _GEN_146 : L0Memory_17; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_247 = count >= 10'h1 & count <= _T_27 ? _GEN_147 : L0Memory_18; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_248 = count >= 10'h1 & count <= _T_27 ? _GEN_148 : L0Memory_19; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_249 = count >= 10'h1 & count <= _T_27 ? _GEN_149 : L0Memory_20; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_250 = count >= 10'h1 & count <= _T_27 ? _GEN_150 : L0Memory_21; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_251 = count >= 10'h1 & count <= _T_27 ? _GEN_151 : L0Memory_22; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_252 = count >= 10'h1 & count <= _T_27 ? _GEN_152 : L0Memory_23; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_253 = count >= 10'h1 & count <= _T_27 ? _GEN_153 : L0Memory_24; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_254 = count >= 10'h1 & count <= _T_27 ? _GEN_154 : L0Memory_25; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_255 = count >= 10'h1 & count <= _T_27 ? _GEN_155 : L0Memory_26; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_256 = count >= 10'h1 & count <= _T_27 ? _GEN_156 : L0Memory_27; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_257 = count >= 10'h1 & count <= _T_27 ? _GEN_157 : L0Memory_28; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_258 = count >= 10'h1 & count <= _T_27 ? _GEN_158 : L0Memory_29; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_259 = count >= 10'h1 & count <= _T_27 ? _GEN_159 : L0Memory_30; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_260 = count >= 10'h1 & count <= _T_27 ? _GEN_160 : L0Memory_31; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_261 = count >= 10'h1 & count <= _T_27 ? _GEN_161 : L0Memory_32; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_262 = count >= 10'h1 & count <= _T_27 ? _GEN_162 : L0Memory_33; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_263 = count >= 10'h1 & count <= _T_27 ? _GEN_163 : L0Memory_34; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_264 = count >= 10'h1 & count <= _T_27 ? _GEN_164 : L0Memory_35; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_265 = count >= 10'h1 & count <= _T_27 ? _GEN_165 : L0Memory_36; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_266 = count >= 10'h1 & count <= _T_27 ? _GEN_166 : L0Memory_37; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_267 = count >= 10'h1 & count <= _T_27 ? _GEN_167 : L0Memory_38; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_268 = count >= 10'h1 & count <= _T_27 ? _GEN_168 : L0Memory_39; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_269 = count >= 10'h1 & count <= _T_27 ? _GEN_169 : L0Memory_40; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_270 = count >= 10'h1 & count <= _T_27 ? _GEN_170 : L0Memory_41; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_271 = count >= 10'h1 & count <= _T_27 ? _GEN_171 : L0Memory_42; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_272 = count >= 10'h1 & count <= _T_27 ? _GEN_172 : L0Memory_43; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_273 = count >= 10'h1 & count <= _T_27 ? _GEN_173 : L0Memory_44; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_274 = count >= 10'h1 & count <= _T_27 ? _GEN_174 : L0Memory_45; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_275 = count >= 10'h1 & count <= _T_27 ? _GEN_175 : L0Memory_46; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_276 = count >= 10'h1 & count <= _T_27 ? _GEN_176 : L0Memory_47; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_277 = count >= 10'h1 & count <= _T_27 ? _GEN_177 : L0Memory_48; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_278 = count >= 10'h1 & count <= _T_27 ? _GEN_178 : L0Memory_49; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_279 = count >= 10'h1 & count <= _T_27 ? _GEN_179 : L0Memory_50; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_280 = count >= 10'h1 & count <= _T_27 ? _GEN_180 : L0Memory_51; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_281 = count >= 10'h1 & count <= _T_27 ? _GEN_181 : L0Memory_52; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_282 = count >= 10'h1 & count <= _T_27 ? _GEN_182 : L0Memory_53; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_283 = count >= 10'h1 & count <= _T_27 ? _GEN_183 : L0Memory_54; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_284 = count >= 10'h1 & count <= _T_27 ? _GEN_184 : L0Memory_55; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_285 = count >= 10'h1 & count <= _T_27 ? _GEN_185 : L0Memory_56; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_286 = count >= 10'h1 & count <= _T_27 ? _GEN_186 : L0Memory_57; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_287 = count >= 10'h1 & count <= _T_27 ? _GEN_187 : L0Memory_58; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_288 = count >= 10'h1 & count <= _T_27 ? _GEN_188 : L0Memory_59; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_289 = count >= 10'h1 & count <= _T_27 ? _GEN_189 : L0Memory_60; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_290 = count >= 10'h1 & count <= _T_27 ? _GEN_190 : L0Memory_61; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_291 = count >= 10'h1 & count <= _T_27 ? _GEN_191 : L0Memory_62; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_292 = count >= 10'h1 & count <= _T_27 ? _GEN_192 : L0Memory_63; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_293 = count >= 10'h1 & count <= _T_27 ? _GEN_193 : L0Memory_64; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_294 = count >= 10'h1 & count <= _T_27 ? _GEN_194 : L0Memory_65; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_295 = count >= 10'h1 & count <= _T_27 ? _GEN_195 : L0Memory_66; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_296 = count >= 10'h1 & count <= _T_27 ? _GEN_196 : L0Memory_67; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_297 = count >= 10'h1 & count <= _T_27 ? _GEN_197 : L0Memory_68; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_298 = count >= 10'h1 & count <= _T_27 ? _GEN_198 : L0Memory_69; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_299 = count >= 10'h1 & count <= _T_27 ? _GEN_199 : L0Memory_70; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_300 = count >= 10'h1 & count <= _T_27 ? _GEN_200 : L0Memory_71; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_301 = count >= 10'h1 & count <= _T_27 ? _GEN_201 : L0Memory_72; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_302 = count >= 10'h1 & count <= _T_27 ? _GEN_202 : L0Memory_73; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_303 = count >= 10'h1 & count <= _T_27 ? _GEN_203 : L0Memory_74; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_304 = count >= 10'h1 & count <= _T_27 ? _GEN_204 : L0Memory_75; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_305 = count >= 10'h1 & count <= _T_27 ? _GEN_205 : L0Memory_76; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_306 = count >= 10'h1 & count <= _T_27 ? _GEN_206 : L0Memory_77; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_307 = count >= 10'h1 & count <= _T_27 ? _GEN_207 : L0Memory_78; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_308 = count >= 10'h1 & count <= _T_27 ? _GEN_208 : L0Memory_79; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_309 = count >= 10'h1 & count <= _T_27 ? _GEN_209 : L0Memory_80; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_310 = count >= 10'h1 & count <= _T_27 ? _GEN_210 : L0Memory_81; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_311 = count >= 10'h1 & count <= _T_27 ? _GEN_211 : L0Memory_82; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_312 = count >= 10'h1 & count <= _T_27 ? _GEN_212 : L0Memory_83; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_313 = count >= 10'h1 & count <= _T_27 ? _GEN_213 : L0Memory_84; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_314 = count >= 10'h1 & count <= _T_27 ? _GEN_214 : L0Memory_85; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_315 = count >= 10'h1 & count <= _T_27 ? _GEN_215 : L0Memory_86; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_316 = count >= 10'h1 & count <= _T_27 ? _GEN_216 : L0Memory_87; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_317 = count >= 10'h1 & count <= _T_27 ? _GEN_217 : L0Memory_88; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_318 = count >= 10'h1 & count <= _T_27 ? _GEN_218 : L0Memory_89; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_319 = count >= 10'h1 & count <= _T_27 ? _GEN_219 : L0Memory_90; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_320 = count >= 10'h1 & count <= _T_27 ? _GEN_220 : L0Memory_91; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_321 = count >= 10'h1 & count <= _T_27 ? _GEN_221 : L0Memory_92; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_322 = count >= 10'h1 & count <= _T_27 ? _GEN_222 : L0Memory_93; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_323 = count >= 10'h1 & count <= _T_27 ? _GEN_223 : L0Memory_94; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_324 = count >= 10'h1 & count <= _T_27 ? _GEN_224 : L0Memory_95; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_325 = count >= 10'h1 & count <= _T_27 ? _GEN_225 : L0Memory_96; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_326 = count >= 10'h1 & count <= _T_27 ? _GEN_226 : L0Memory_97; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_327 = count >= 10'h1 & count <= _T_27 ? _GEN_227 : L0Memory_98; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_328 = count >= 10'h1 & count <= _T_27 ? _GEN_228 : L0Memory_99; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [5:0] _GEN_329 = count >= 10'h1 & count <= _T_27 ? _L0Index_T_2 : _GEN_128; // @[PEArray.scala 198:59 PEArray.scala 200:17]
  wire [9:0] _GEN_330 = _T_24 ? 10'h0 : _GEN_127; // @[PEArray.scala 202:32 PEArray.scala 203:15]
  wire [2:0] _GEN_331 = _T_24 ? 3'h0 : state; // @[PEArray.scala 202:32 PEArray.scala 204:15 PEArray.scala 100:22]
  wire [9:0] _GEN_865 = {{4'd0}, GRU_out_width}; // @[PEArray.scala 220:19]
  wire [9:0] _GEN_0 = count % _GEN_865; // @[PEArray.scala 220:19]
  wire [5:0] _T_36 = _GEN_0[5:0]; // @[PEArray.scala 220:19]
  wire [5:0] _T_38 = GRU_out_width - 6'h1; // @[PEArray.scala 220:55]
  wire [5:0] _GEN_334 = _T_36 == _T_38 ? _L0Index_T_2 : 6'h0; // @[PEArray.scala 220:62 PEArray.scala 221:17 PEArray.scala 214:15]
  wire [5:0] _GEN_346 = _T_41 ? _GEN_334 : L0Index; // @[Conditional.scala 39:67 PEArray.scala 39:24]
  wire [9:0] _GEN_347 = _T_41 ? _GEN_330 : count; // @[Conditional.scala 39:67 PEArray.scala 101:22]
  wire [2:0] _GEN_348 = _T_41 ? _GEN_331 : state; // @[Conditional.scala 39:67 PEArray.scala 100:22]
  wire [5:0] _GEN_353 = _T_31 ? _GEN_334 : _GEN_346; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_354 = _T_31 ? _GEN_330 : _GEN_347; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_355 = _T_31 ? _GEN_331 : _GEN_348; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_356 = _T_22 ? _GEN_330 : _GEN_354; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_357 = _T_22 ? _GEN_329 : _GEN_353; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_458 = _T_22 ? _GEN_331 : _GEN_355; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_690 = _T_3 ? _GEN_118 : {{2'd0}, GRU_out_width}; // @[Conditional.scala 40:58 PEArray.scala 104:26]
  FP16MulAdder FP16MAC ( // @[PEArray.scala 72:23]
    .io_a(FP16MAC_io_a),
    .io_b(FP16MAC_io_b),
    .io_c(FP16MAC_io_c),
    .io_out(FP16MAC_io_out)
  );
  assign io_ToRightPE = mux3out_reg; // @[PEArray.scala 95:16]
  assign io_ToBelowPE = mux2out_reg; // @[PEArray.scala 94:16]
  assign FP16MAC_io_a = sel1 ? io_FromL1 : io_FromLeftPE; // @[PEArray.scala 50:14 PEArray.scala 50:23 PEArray.scala 51:24]
  assign FP16MAC_io_b = sel5 ? mux4out : _GEN_105; // @[PEArray.scala 77:13 PEArray.scala 78:18 PEArray.scala 81:18]
  assign FP16MAC_io_c = sel5 ? _GEN_105 : mux4out; // @[PEArray.scala 77:13 PEArray.scala 79:18 PEArray.scala 82:18]
  always @(posedge clock) begin
    if (reset) begin // @[PEArray.scala 39:24]
      L0Index <= 6'h0; // @[PEArray.scala 39:24]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h1; // @[PEArray.scala 159:15]
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h6; // @[PEArray.scala 181:15]
      end else begin
        L0Index <= _GEN_357;
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_0 <= _GEN_229;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_1 <= _GEN_230;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_2 <= _GEN_231;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_3 <= _GEN_232;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_4 <= _GEN_233;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_5 <= _GEN_234;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_6 <= _GEN_235;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_7 <= _GEN_236;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_8 <= _GEN_237;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_9 <= _GEN_238;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_10 <= _GEN_239;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_11 <= _GEN_240;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_12 <= _GEN_241;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_13 <= _GEN_242;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_14 <= _GEN_243;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_15 <= _GEN_244;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_16 <= _GEN_245;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_17 <= _GEN_246;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_18 <= _GEN_247;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_19 <= _GEN_248;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_20 <= _GEN_249;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_21 <= _GEN_250;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_22 <= _GEN_251;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_23 <= _GEN_252;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_24 <= _GEN_253;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_25 <= _GEN_254;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_26 <= _GEN_255;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_27 <= _GEN_256;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_28 <= _GEN_257;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_29 <= _GEN_258;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_30 <= _GEN_259;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_31 <= _GEN_260;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_32 <= _GEN_261;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_33 <= _GEN_262;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_34 <= _GEN_263;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_35 <= _GEN_264;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_36 <= _GEN_265;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_37 <= _GEN_266;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_38 <= _GEN_267;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_39 <= _GEN_268;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_40 <= _GEN_269;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_41 <= _GEN_270;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_42 <= _GEN_271;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_43 <= _GEN_272;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_44 <= _GEN_273;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_45 <= _GEN_274;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_46 <= _GEN_275;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_47 <= _GEN_276;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_48 <= _GEN_277;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_49 <= _GEN_278;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_50 <= _GEN_279;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_51 <= _GEN_280;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_52 <= _GEN_281;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_53 <= _GEN_282;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_54 <= _GEN_283;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_55 <= _GEN_284;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_56 <= _GEN_285;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_57 <= _GEN_286;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_58 <= _GEN_287;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_59 <= _GEN_288;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_60 <= _GEN_289;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_61 <= _GEN_290;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_62 <= _GEN_291;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_63 <= _GEN_292;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_64 <= _GEN_293;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_65 <= _GEN_294;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_66 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_67 <= _GEN_296;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_68 <= _GEN_297;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_69 <= _GEN_298;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_70 <= _GEN_299;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_71 <= _GEN_300;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_72 <= _GEN_301;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_73 <= _GEN_302;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_74 <= _GEN_303;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_75 <= _GEN_304;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_76 <= _GEN_305;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_77 <= _GEN_306;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_78 <= _GEN_307;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_79 <= _GEN_308;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_80 <= _GEN_309;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_81 <= _GEN_310;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_82 <= _GEN_311;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_83 <= _GEN_312;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_84 <= _GEN_313;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_85 <= _GEN_314;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_86 <= _GEN_315;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_87 <= _GEN_316;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_88 <= _GEN_317;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_89 <= _GEN_318;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_90 <= _GEN_319;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_91 <= _GEN_320;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_92 <= _GEN_321;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_93 <= _GEN_322;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_94 <= _GEN_323;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_95 <= _GEN_324;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_96 <= _GEN_325;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_97 <= _GEN_326;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_98 <= _GEN_327;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_99 <= _GEN_328;
          end
        end
      end
    end
    if (reset) begin // @[PEArray.scala 100:22]
      state <= 3'h0; // @[PEArray.scala 100:22]
    end else if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[8]) begin // @[PEArray.scala 116:57]
        state <= 3'h1;
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      if (count == 10'h33) begin // @[PEArray.scala 164:27]
        state <= 3'h0; // @[PEArray.scala 166:15]
      end
    end else if (_T_16) begin // @[Conditional.scala 39:67]
      state <= _GEN_126;
    end else begin
      state <= _GEN_458;
    end
    if (reset) begin // @[PEArray.scala 90:28]
      mux2out_reg <= 16'h0; // @[PEArray.scala 90:28]
    end else begin
      mux2out_reg <= MAC_out; // @[PEArray.scala 90:28]
    end
    if (reset) begin // @[PEArray.scala 91:28]
      mux3out_reg <= 16'h0; // @[PEArray.scala 91:28]
    end else if (sel3) begin // @[PEArray.scala 56:14]
      mux3out_reg <= MAC_out; // @[PEArray.scala 56:23]
    end else if (sel1) begin // @[PEArray.scala 50:14]
      mux3out_reg <= io_FromL1; // @[PEArray.scala 50:23]
    end else begin
      mux3out_reg <= io_FromLeftPE; // @[PEArray.scala 51:24]
    end
    if (reset) begin // @[PEArray.scala 101:22]
      count <= 10'h0; // @[PEArray.scala 101:22]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        if (count == 10'h33) begin // @[PEArray.scala 164:27]
          count <= 10'h0; // @[PEArray.scala 165:15]
        end else begin
          count <= _GEN_120;
        end
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        count <= _GEN_125;
      end else begin
        count <= _GEN_356;
      end
    end
    GRU_out_width <= _GEN_690[5:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  L0Index = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  L0Memory_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  L0Memory_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  L0Memory_2 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  L0Memory_3 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  L0Memory_4 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  L0Memory_5 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  L0Memory_6 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  L0Memory_7 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  L0Memory_8 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  L0Memory_9 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  L0Memory_10 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  L0Memory_11 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  L0Memory_12 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  L0Memory_13 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  L0Memory_14 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  L0Memory_15 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  L0Memory_16 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  L0Memory_17 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  L0Memory_18 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  L0Memory_19 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  L0Memory_20 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  L0Memory_21 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  L0Memory_22 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  L0Memory_23 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  L0Memory_24 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  L0Memory_25 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  L0Memory_26 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  L0Memory_27 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  L0Memory_28 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  L0Memory_29 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  L0Memory_30 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  L0Memory_31 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  L0Memory_32 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  L0Memory_33 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  L0Memory_34 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  L0Memory_35 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  L0Memory_36 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  L0Memory_37 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  L0Memory_38 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  L0Memory_39 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  L0Memory_40 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  L0Memory_41 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  L0Memory_42 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  L0Memory_43 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  L0Memory_44 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  L0Memory_45 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  L0Memory_46 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  L0Memory_47 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  L0Memory_48 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  L0Memory_49 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  L0Memory_50 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  L0Memory_51 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  L0Memory_52 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  L0Memory_53 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  L0Memory_54 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  L0Memory_55 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  L0Memory_56 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  L0Memory_57 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  L0Memory_58 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  L0Memory_59 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  L0Memory_60 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  L0Memory_61 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  L0Memory_62 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  L0Memory_63 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  L0Memory_64 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  L0Memory_65 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  L0Memory_66 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  L0Memory_67 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  L0Memory_68 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  L0Memory_69 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  L0Memory_70 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  L0Memory_71 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  L0Memory_72 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  L0Memory_73 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  L0Memory_74 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  L0Memory_75 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  L0Memory_76 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  L0Memory_77 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  L0Memory_78 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  L0Memory_79 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  L0Memory_80 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  L0Memory_81 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  L0Memory_82 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  L0Memory_83 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  L0Memory_84 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  L0Memory_85 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  L0Memory_86 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  L0Memory_87 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  L0Memory_88 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  L0Memory_89 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  L0Memory_90 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  L0Memory_91 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  L0Memory_92 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  L0Memory_93 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  L0Memory_94 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  L0Memory_95 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  L0Memory_96 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  L0Memory_97 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  L0Memory_98 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  L0Memory_99 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  state = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  mux2out_reg = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  mux3out_reg = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  count = _RAND_104[9:0];
  _RAND_105 = {1{`RANDOM}};
  GRU_out_width = _RAND_105[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PE_11(
  input         clock,
  input         reset,
  input  [15:0] io_FromAbovePE,
  input  [15:0] io_FromLeftPE,
  input  [15:0] io_FromL1,
  input  [2:0]  io_control_signal_control,
  input  [9:0]  io_control_signal_count,
  input  [5:0]  io_control_signal_L0index,
  input  [11:0] io_control_signal_mask,
  input  [7:0]  io_control_signal_gru_out_width,
  output [15:0] io_ToRightPE,
  output [15:0] io_ToBelowPE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] FP16MAC_io_a; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_b; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_c; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_out; // @[PEArray.scala 72:23]
  reg [5:0] L0Index; // @[PEArray.scala 39:24]
  reg [15:0] L0Memory_0; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_1; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_2; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_3; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_4; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_5; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_6; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_7; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_8; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_9; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_10; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_11; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_12; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_13; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_14; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_15; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_16; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_17; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_18; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_19; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_20; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_21; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_22; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_23; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_24; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_25; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_26; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_27; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_28; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_29; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_30; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_31; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_32; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_33; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_34; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_35; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_36; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_37; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_38; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_39; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_40; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_41; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_42; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_43; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_44; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_45; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_46; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_47; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_48; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_49; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_50; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_51; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_52; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_53; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_54; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_55; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_56; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_57; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_58; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_59; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_60; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_61; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_62; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_63; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_64; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_65; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_66; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_67; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_68; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_69; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_70; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_71; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_72; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_73; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_74; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_75; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_76; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_77; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_78; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_79; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_80; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_81; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_82; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_83; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_84; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_85; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_86; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_87; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_88; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_89; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_90; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_91; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_92; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_93; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_94; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_95; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_96; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_97; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_98; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_99; // @[PEArray.scala 40:21]
  reg [2:0] state; // @[PEArray.scala 100:22]
  wire  _T_3 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_12 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_16 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_22 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_31 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_41 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_342 = _T_41 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 231:12 PEArray.scala 32:8]
  wire  _GEN_349 = _T_31 ? 1'h0 : _GEN_342; // @[Conditional.scala 39:67 PEArray.scala 208:12]
  wire  _GEN_459 = _T_22 | _GEN_349; // @[Conditional.scala 39:67 PEArray.scala 32:8]
  wire  _GEN_463 = _T_16 ? 1'h0 : _GEN_459; // @[Conditional.scala 39:67]
  wire  _GEN_572 = _T_12 | _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 149:12]
  wire  sel1 = _T_3 | _GEN_572; // @[Conditional.scala 40:58 PEArray.scala 108:12]
  wire [15:0] MAC_out = FP16MAC_io_out; // @[PEArray.scala 47:21 PEArray.scala 85:11]
  wire  _GEN_465 = _T_16 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 177:12]
  wire  _GEN_580 = _T_12 | _GEN_465; // @[Conditional.scala 39:67 PEArray.scala 34:8]
  wire  sel3 = _T_3 | _GEN_580; // @[Conditional.scala 40:58 PEArray.scala 110:12]
  wire [1:0] _GEN_344 = _T_41 ? 2'h2 : 2'h0; // @[Conditional.scala 39:67 PEArray.scala 233:12 PEArray.scala 35:8]
  wire [1:0] _GEN_351 = _T_31 ? 2'h2 : _GEN_344; // @[Conditional.scala 39:67 PEArray.scala 210:12]
  wire [1:0] _GEN_461 = _T_22 ? 2'h0 : _GEN_351; // @[Conditional.scala 39:67 PEArray.scala 35:8]
  wire [1:0] _GEN_466 = _T_16 ? 2'h0 : _GEN_461; // @[Conditional.scala 39:67 PEArray.scala 178:12]
  wire [1:0] _GEN_574 = _T_12 ? 2'h1 : _GEN_466; // @[Conditional.scala 39:67]
  wire [1:0] sel4 = _T_3 ? 2'h0 : _GEN_574; // @[Conditional.scala 40:58 PEArray.scala 111:12]
  wire [15:0] _GEN_3 = sel4 == 2'h2 ? io_FromL1 : 16'h0; // @[PEArray.scala 65:28 PEArray.scala 66:15 PEArray.scala 69:15]
  wire [15:0] _GEN_4 = sel4 == 2'h1 ? io_FromAbovePE : _GEN_3; // @[PEArray.scala 62:28 PEArray.scala 63:15]
  wire [15:0] mux4out = sel4 == 2'h0 ? 16'h0 : _GEN_4; // @[PEArray.scala 59:22 PEArray.scala 60:13]
  wire [15:0] _GEN_7 = 6'h1 == L0Index ? L0Memory_1 : L0Memory_0; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_8 = 6'h2 == L0Index ? L0Memory_2 : _GEN_7; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_9 = 6'h3 == L0Index ? L0Memory_3 : _GEN_8; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_10 = 6'h4 == L0Index ? L0Memory_4 : _GEN_9; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_11 = 6'h5 == L0Index ? L0Memory_5 : _GEN_10; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_12 = 6'h6 == L0Index ? L0Memory_6 : _GEN_11; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_13 = 6'h7 == L0Index ? L0Memory_7 : _GEN_12; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_14 = 6'h8 == L0Index ? L0Memory_8 : _GEN_13; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_15 = 6'h9 == L0Index ? L0Memory_9 : _GEN_14; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_16 = 6'ha == L0Index ? L0Memory_10 : _GEN_15; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_17 = 6'hb == L0Index ? L0Memory_11 : _GEN_16; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_18 = 6'hc == L0Index ? L0Memory_12 : _GEN_17; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_19 = 6'hd == L0Index ? L0Memory_13 : _GEN_18; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_20 = 6'he == L0Index ? L0Memory_14 : _GEN_19; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_21 = 6'hf == L0Index ? L0Memory_15 : _GEN_20; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_22 = 6'h10 == L0Index ? L0Memory_16 : _GEN_21; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_23 = 6'h11 == L0Index ? L0Memory_17 : _GEN_22; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_24 = 6'h12 == L0Index ? L0Memory_18 : _GEN_23; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_25 = 6'h13 == L0Index ? L0Memory_19 : _GEN_24; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_26 = 6'h14 == L0Index ? L0Memory_20 : _GEN_25; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_27 = 6'h15 == L0Index ? L0Memory_21 : _GEN_26; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_28 = 6'h16 == L0Index ? L0Memory_22 : _GEN_27; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_29 = 6'h17 == L0Index ? L0Memory_23 : _GEN_28; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_30 = 6'h18 == L0Index ? L0Memory_24 : _GEN_29; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_31 = 6'h19 == L0Index ? L0Memory_25 : _GEN_30; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_32 = 6'h1a == L0Index ? L0Memory_26 : _GEN_31; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_33 = 6'h1b == L0Index ? L0Memory_27 : _GEN_32; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_34 = 6'h1c == L0Index ? L0Memory_28 : _GEN_33; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_35 = 6'h1d == L0Index ? L0Memory_29 : _GEN_34; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_36 = 6'h1e == L0Index ? L0Memory_30 : _GEN_35; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_37 = 6'h1f == L0Index ? L0Memory_31 : _GEN_36; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_38 = 6'h20 == L0Index ? L0Memory_32 : _GEN_37; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_39 = 6'h21 == L0Index ? L0Memory_33 : _GEN_38; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_40 = 6'h22 == L0Index ? L0Memory_34 : _GEN_39; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_41 = 6'h23 == L0Index ? L0Memory_35 : _GEN_40; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_42 = 6'h24 == L0Index ? L0Memory_36 : _GEN_41; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_43 = 6'h25 == L0Index ? L0Memory_37 : _GEN_42; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_44 = 6'h26 == L0Index ? L0Memory_38 : _GEN_43; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_45 = 6'h27 == L0Index ? L0Memory_39 : _GEN_44; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_46 = 6'h28 == L0Index ? L0Memory_40 : _GEN_45; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_47 = 6'h29 == L0Index ? L0Memory_41 : _GEN_46; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_48 = 6'h2a == L0Index ? L0Memory_42 : _GEN_47; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_49 = 6'h2b == L0Index ? L0Memory_43 : _GEN_48; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_50 = 6'h2c == L0Index ? L0Memory_44 : _GEN_49; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_51 = 6'h2d == L0Index ? L0Memory_45 : _GEN_50; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_52 = 6'h2e == L0Index ? L0Memory_46 : _GEN_51; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_53 = 6'h2f == L0Index ? L0Memory_47 : _GEN_52; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_54 = 6'h30 == L0Index ? L0Memory_48 : _GEN_53; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_55 = 6'h31 == L0Index ? L0Memory_49 : _GEN_54; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_56 = 6'h32 == L0Index ? L0Memory_50 : _GEN_55; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_57 = 6'h33 == L0Index ? L0Memory_51 : _GEN_56; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_58 = 6'h34 == L0Index ? L0Memory_52 : _GEN_57; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_59 = 6'h35 == L0Index ? L0Memory_53 : _GEN_58; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_60 = 6'h36 == L0Index ? L0Memory_54 : _GEN_59; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_61 = 6'h37 == L0Index ? L0Memory_55 : _GEN_60; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_62 = 6'h38 == L0Index ? L0Memory_56 : _GEN_61; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_63 = 6'h39 == L0Index ? L0Memory_57 : _GEN_62; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_64 = 6'h3a == L0Index ? L0Memory_58 : _GEN_63; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_65 = 6'h3b == L0Index ? L0Memory_59 : _GEN_64; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_66 = 6'h3c == L0Index ? L0Memory_60 : _GEN_65; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_67 = 6'h3d == L0Index ? L0Memory_61 : _GEN_66; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_68 = 6'h3e == L0Index ? L0Memory_62 : _GEN_67; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_69 = 6'h3f == L0Index ? L0Memory_63 : _GEN_68; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [6:0] _GEN_793 = {{1'd0}, L0Index}; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_70 = 7'h40 == _GEN_793 ? L0Memory_64 : _GEN_69; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_71 = 7'h41 == _GEN_793 ? L0Memory_65 : _GEN_70; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_72 = 7'h42 == _GEN_793 ? L0Memory_66 : _GEN_71; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_73 = 7'h43 == _GEN_793 ? L0Memory_67 : _GEN_72; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_74 = 7'h44 == _GEN_793 ? L0Memory_68 : _GEN_73; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_75 = 7'h45 == _GEN_793 ? L0Memory_69 : _GEN_74; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_76 = 7'h46 == _GEN_793 ? L0Memory_70 : _GEN_75; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_77 = 7'h47 == _GEN_793 ? L0Memory_71 : _GEN_76; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_78 = 7'h48 == _GEN_793 ? L0Memory_72 : _GEN_77; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_79 = 7'h49 == _GEN_793 ? L0Memory_73 : _GEN_78; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_80 = 7'h4a == _GEN_793 ? L0Memory_74 : _GEN_79; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_81 = 7'h4b == _GEN_793 ? L0Memory_75 : _GEN_80; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_82 = 7'h4c == _GEN_793 ? L0Memory_76 : _GEN_81; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_83 = 7'h4d == _GEN_793 ? L0Memory_77 : _GEN_82; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_84 = 7'h4e == _GEN_793 ? L0Memory_78 : _GEN_83; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_85 = 7'h4f == _GEN_793 ? L0Memory_79 : _GEN_84; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_86 = 7'h50 == _GEN_793 ? L0Memory_80 : _GEN_85; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_87 = 7'h51 == _GEN_793 ? L0Memory_81 : _GEN_86; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_88 = 7'h52 == _GEN_793 ? L0Memory_82 : _GEN_87; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_89 = 7'h53 == _GEN_793 ? L0Memory_83 : _GEN_88; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_90 = 7'h54 == _GEN_793 ? L0Memory_84 : _GEN_89; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_91 = 7'h55 == _GEN_793 ? L0Memory_85 : _GEN_90; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_92 = 7'h56 == _GEN_793 ? L0Memory_86 : _GEN_91; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_93 = 7'h57 == _GEN_793 ? L0Memory_87 : _GEN_92; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_94 = 7'h58 == _GEN_793 ? L0Memory_88 : _GEN_93; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_95 = 7'h59 == _GEN_793 ? L0Memory_89 : _GEN_94; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_96 = 7'h5a == _GEN_793 ? L0Memory_90 : _GEN_95; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_97 = 7'h5b == _GEN_793 ? L0Memory_91 : _GEN_96; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_98 = 7'h5c == _GEN_793 ? L0Memory_92 : _GEN_97; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_99 = 7'h5d == _GEN_793 ? L0Memory_93 : _GEN_98; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_100 = 7'h5e == _GEN_793 ? L0Memory_94 : _GEN_99; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_101 = 7'h5f == _GEN_793 ? L0Memory_95 : _GEN_100; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_102 = 7'h60 == _GEN_793 ? L0Memory_96 : _GEN_101; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_103 = 7'h61 == _GEN_793 ? L0Memory_97 : _GEN_102; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_104 = 7'h62 == _GEN_793 ? L0Memory_98 : _GEN_103; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_105 = 7'h63 == _GEN_793 ? L0Memory_99 : _GEN_104; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire  _GEN_575 = _T_12 ? 1'h0 : _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 157:12]
  wire  sel5 = _T_3 ? 1'h0 : _GEN_575; // @[Conditional.scala 40:58 PEArray.scala 112:12]
  reg [15:0] mux2out_reg; // @[PEArray.scala 90:28]
  reg [15:0] mux3out_reg; // @[PEArray.scala 91:28]
  reg [9:0] count; // @[PEArray.scala 101:22]
  reg [9:0] count_max; // @[PEArray.scala 102:22]
  reg [5:0] L0index_begin; // @[PEArray.scala 103:26]
  reg [5:0] GRU_out_width; // @[PEArray.scala 104:26]
  wire  _T_6 = 3'h0 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_7 = 3'h1 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_8 = 3'h2 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_9 = 3'h3 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_10 = 3'h4 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_11 = 3'h5 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_109 = _T_11 ? 3'h5 : state; // @[Conditional.scala 39:67 PEArray.scala 140:19 PEArray.scala 100:22]
  wire [2:0] _GEN_110 = _T_10 ? 3'h4 : _GEN_109; // @[Conditional.scala 39:67 PEArray.scala 136:19]
  wire [2:0] _GEN_111 = _T_9 ? 3'h3 : _GEN_110; // @[Conditional.scala 39:67 PEArray.scala 132:19]
  wire [2:0] _GEN_112 = _T_8 ? 3'h2 : _GEN_111; // @[Conditional.scala 39:67 PEArray.scala 128:19]
  wire [2:0] _GEN_113 = _T_7 ? 3'h1 : _GEN_112; // @[Conditional.scala 39:67 PEArray.scala 124:19]
  wire [7:0] _GEN_118 = io_control_signal_mask[8] ? io_control_signal_gru_out_width : {{2'd0}, GRU_out_width}; // @[PEArray.scala 116:57 PEArray.scala 145:23 PEArray.scala 104:26]
  wire [9:0] _count_T_1 = count + 10'h1; // @[PEArray.scala 162:24]
  wire [9:0] _GEN_120 = count != 10'h33 ? _count_T_1 : count; // @[PEArray.scala 161:27 PEArray.scala 162:15 PEArray.scala 101:22]
  wire [9:0] _GEN_124 = count != 10'h188 ? _count_T_1 : count; // @[PEArray.scala 183:28 PEArray.scala 184:15 PEArray.scala 101:22]
  wire [9:0] _GEN_125 = count == 10'h188 ? 10'h0 : _GEN_124; // @[PEArray.scala 186:28 PEArray.scala 187:15]
  wire [2:0] _GEN_126 = count == 10'h188 ? 3'h0 : state; // @[PEArray.scala 186:28 PEArray.scala 188:15 PEArray.scala 100:22]
  wire [9:0] _GEN_127 = count != count_max ? _count_T_1 : count; // @[PEArray.scala 192:32 PEArray.scala 193:15 PEArray.scala 101:22]
  wire [5:0] _GEN_128 = count == 10'h0 ? L0index_begin : L0Index; // @[PEArray.scala 195:26 PEArray.scala 196:17 PEArray.scala 39:24]
  wire [9:0] _T_27 = count_max - 10'h1; // @[PEArray.scala 198:51]
  wire [15:0] _GEN_129 = 6'h0 == L0Index ? io_FromL1 : L0Memory_0; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_130 = 6'h1 == L0Index ? io_FromL1 : L0Memory_1; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_131 = 6'h2 == L0Index ? io_FromL1 : L0Memory_2; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_132 = 6'h3 == L0Index ? io_FromL1 : L0Memory_3; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_133 = 6'h4 == L0Index ? io_FromL1 : L0Memory_4; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_134 = 6'h5 == L0Index ? io_FromL1 : L0Memory_5; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_135 = 6'h6 == L0Index ? io_FromL1 : L0Memory_6; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_136 = 6'h7 == L0Index ? io_FromL1 : L0Memory_7; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_137 = 6'h8 == L0Index ? io_FromL1 : L0Memory_8; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_138 = 6'h9 == L0Index ? io_FromL1 : L0Memory_9; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_139 = 6'ha == L0Index ? io_FromL1 : L0Memory_10; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_140 = 6'hb == L0Index ? io_FromL1 : L0Memory_11; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_141 = 6'hc == L0Index ? io_FromL1 : L0Memory_12; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_142 = 6'hd == L0Index ? io_FromL1 : L0Memory_13; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_143 = 6'he == L0Index ? io_FromL1 : L0Memory_14; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_144 = 6'hf == L0Index ? io_FromL1 : L0Memory_15; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_145 = 6'h10 == L0Index ? io_FromL1 : L0Memory_16; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_146 = 6'h11 == L0Index ? io_FromL1 : L0Memory_17; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_147 = 6'h12 == L0Index ? io_FromL1 : L0Memory_18; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_148 = 6'h13 == L0Index ? io_FromL1 : L0Memory_19; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_149 = 6'h14 == L0Index ? io_FromL1 : L0Memory_20; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_150 = 6'h15 == L0Index ? io_FromL1 : L0Memory_21; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_151 = 6'h16 == L0Index ? io_FromL1 : L0Memory_22; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_152 = 6'h17 == L0Index ? io_FromL1 : L0Memory_23; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_153 = 6'h18 == L0Index ? io_FromL1 : L0Memory_24; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_154 = 6'h19 == L0Index ? io_FromL1 : L0Memory_25; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_155 = 6'h1a == L0Index ? io_FromL1 : L0Memory_26; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_156 = 6'h1b == L0Index ? io_FromL1 : L0Memory_27; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_157 = 6'h1c == L0Index ? io_FromL1 : L0Memory_28; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_158 = 6'h1d == L0Index ? io_FromL1 : L0Memory_29; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_159 = 6'h1e == L0Index ? io_FromL1 : L0Memory_30; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_160 = 6'h1f == L0Index ? io_FromL1 : L0Memory_31; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_161 = 6'h20 == L0Index ? io_FromL1 : L0Memory_32; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_162 = 6'h21 == L0Index ? io_FromL1 : L0Memory_33; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_163 = 6'h22 == L0Index ? io_FromL1 : L0Memory_34; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_164 = 6'h23 == L0Index ? io_FromL1 : L0Memory_35; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_165 = 6'h24 == L0Index ? io_FromL1 : L0Memory_36; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_166 = 6'h25 == L0Index ? io_FromL1 : L0Memory_37; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_167 = 6'h26 == L0Index ? io_FromL1 : L0Memory_38; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_168 = 6'h27 == L0Index ? io_FromL1 : L0Memory_39; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_169 = 6'h28 == L0Index ? io_FromL1 : L0Memory_40; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_170 = 6'h29 == L0Index ? io_FromL1 : L0Memory_41; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_171 = 6'h2a == L0Index ? io_FromL1 : L0Memory_42; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_172 = 6'h2b == L0Index ? io_FromL1 : L0Memory_43; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_173 = 6'h2c == L0Index ? io_FromL1 : L0Memory_44; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_174 = 6'h2d == L0Index ? io_FromL1 : L0Memory_45; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_175 = 6'h2e == L0Index ? io_FromL1 : L0Memory_46; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_176 = 6'h2f == L0Index ? io_FromL1 : L0Memory_47; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_177 = 6'h30 == L0Index ? io_FromL1 : L0Memory_48; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_178 = 6'h31 == L0Index ? io_FromL1 : L0Memory_49; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_179 = 6'h32 == L0Index ? io_FromL1 : L0Memory_50; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_180 = 6'h33 == L0Index ? io_FromL1 : L0Memory_51; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_181 = 6'h34 == L0Index ? io_FromL1 : L0Memory_52; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_182 = 6'h35 == L0Index ? io_FromL1 : L0Memory_53; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_183 = 6'h36 == L0Index ? io_FromL1 : L0Memory_54; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_184 = 6'h37 == L0Index ? io_FromL1 : L0Memory_55; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_185 = 6'h38 == L0Index ? io_FromL1 : L0Memory_56; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_186 = 6'h39 == L0Index ? io_FromL1 : L0Memory_57; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_187 = 6'h3a == L0Index ? io_FromL1 : L0Memory_58; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_188 = 6'h3b == L0Index ? io_FromL1 : L0Memory_59; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_189 = 6'h3c == L0Index ? io_FromL1 : L0Memory_60; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_190 = 6'h3d == L0Index ? io_FromL1 : L0Memory_61; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_191 = 6'h3e == L0Index ? io_FromL1 : L0Memory_62; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_192 = 6'h3f == L0Index ? io_FromL1 : L0Memory_63; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_193 = 7'h40 == _GEN_793 ? io_FromL1 : L0Memory_64; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_194 = 7'h41 == _GEN_793 ? io_FromL1 : L0Memory_65; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_195 = 7'h42 == _GEN_793 ? io_FromL1 : L0Memory_66; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_196 = 7'h43 == _GEN_793 ? io_FromL1 : L0Memory_67; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_197 = 7'h44 == _GEN_793 ? io_FromL1 : L0Memory_68; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_198 = 7'h45 == _GEN_793 ? io_FromL1 : L0Memory_69; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_199 = 7'h46 == _GEN_793 ? io_FromL1 : L0Memory_70; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_200 = 7'h47 == _GEN_793 ? io_FromL1 : L0Memory_71; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_201 = 7'h48 == _GEN_793 ? io_FromL1 : L0Memory_72; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_202 = 7'h49 == _GEN_793 ? io_FromL1 : L0Memory_73; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_203 = 7'h4a == _GEN_793 ? io_FromL1 : L0Memory_74; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_204 = 7'h4b == _GEN_793 ? io_FromL1 : L0Memory_75; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_205 = 7'h4c == _GEN_793 ? io_FromL1 : L0Memory_76; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_206 = 7'h4d == _GEN_793 ? io_FromL1 : L0Memory_77; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_207 = 7'h4e == _GEN_793 ? io_FromL1 : L0Memory_78; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_208 = 7'h4f == _GEN_793 ? io_FromL1 : L0Memory_79; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_209 = 7'h50 == _GEN_793 ? io_FromL1 : L0Memory_80; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_210 = 7'h51 == _GEN_793 ? io_FromL1 : L0Memory_81; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_211 = 7'h52 == _GEN_793 ? io_FromL1 : L0Memory_82; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_212 = 7'h53 == _GEN_793 ? io_FromL1 : L0Memory_83; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_213 = 7'h54 == _GEN_793 ? io_FromL1 : L0Memory_84; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_214 = 7'h55 == _GEN_793 ? io_FromL1 : L0Memory_85; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_215 = 7'h56 == _GEN_793 ? io_FromL1 : L0Memory_86; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_216 = 7'h57 == _GEN_793 ? io_FromL1 : L0Memory_87; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_217 = 7'h58 == _GEN_793 ? io_FromL1 : L0Memory_88; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_218 = 7'h59 == _GEN_793 ? io_FromL1 : L0Memory_89; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_219 = 7'h5a == _GEN_793 ? io_FromL1 : L0Memory_90; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_220 = 7'h5b == _GEN_793 ? io_FromL1 : L0Memory_91; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_221 = 7'h5c == _GEN_793 ? io_FromL1 : L0Memory_92; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_222 = 7'h5d == _GEN_793 ? io_FromL1 : L0Memory_93; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_223 = 7'h5e == _GEN_793 ? io_FromL1 : L0Memory_94; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_224 = 7'h5f == _GEN_793 ? io_FromL1 : L0Memory_95; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_225 = 7'h60 == _GEN_793 ? io_FromL1 : L0Memory_96; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_226 = 7'h61 == _GEN_793 ? io_FromL1 : L0Memory_97; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_227 = 7'h62 == _GEN_793 ? io_FromL1 : L0Memory_98; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_228 = 7'h63 == _GEN_793 ? io_FromL1 : L0Memory_99; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [5:0] _L0Index_T_2 = L0Index + 6'h1; // @[PEArray.scala 200:28]
  wire [15:0] _GEN_229 = count >= 10'h1 & count <= _T_27 ? _GEN_129 : L0Memory_0; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_230 = count >= 10'h1 & count <= _T_27 ? _GEN_130 : L0Memory_1; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_231 = count >= 10'h1 & count <= _T_27 ? _GEN_131 : L0Memory_2; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_232 = count >= 10'h1 & count <= _T_27 ? _GEN_132 : L0Memory_3; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_233 = count >= 10'h1 & count <= _T_27 ? _GEN_133 : L0Memory_4; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_234 = count >= 10'h1 & count <= _T_27 ? _GEN_134 : L0Memory_5; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_235 = count >= 10'h1 & count <= _T_27 ? _GEN_135 : L0Memory_6; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_236 = count >= 10'h1 & count <= _T_27 ? _GEN_136 : L0Memory_7; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_237 = count >= 10'h1 & count <= _T_27 ? _GEN_137 : L0Memory_8; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_238 = count >= 10'h1 & count <= _T_27 ? _GEN_138 : L0Memory_9; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_239 = count >= 10'h1 & count <= _T_27 ? _GEN_139 : L0Memory_10; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_240 = count >= 10'h1 & count <= _T_27 ? _GEN_140 : L0Memory_11; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_241 = count >= 10'h1 & count <= _T_27 ? _GEN_141 : L0Memory_12; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_242 = count >= 10'h1 & count <= _T_27 ? _GEN_142 : L0Memory_13; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_243 = count >= 10'h1 & count <= _T_27 ? _GEN_143 : L0Memory_14; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_244 = count >= 10'h1 & count <= _T_27 ? _GEN_144 : L0Memory_15; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_245 = count >= 10'h1 & count <= _T_27 ? _GEN_145 : L0Memory_16; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_246 = count >= 10'h1 & count <= _T_27 ? _GEN_146 : L0Memory_17; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_247 = count >= 10'h1 & count <= _T_27 ? _GEN_147 : L0Memory_18; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_248 = count >= 10'h1 & count <= _T_27 ? _GEN_148 : L0Memory_19; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_249 = count >= 10'h1 & count <= _T_27 ? _GEN_149 : L0Memory_20; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_250 = count >= 10'h1 & count <= _T_27 ? _GEN_150 : L0Memory_21; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_251 = count >= 10'h1 & count <= _T_27 ? _GEN_151 : L0Memory_22; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_252 = count >= 10'h1 & count <= _T_27 ? _GEN_152 : L0Memory_23; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_253 = count >= 10'h1 & count <= _T_27 ? _GEN_153 : L0Memory_24; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_254 = count >= 10'h1 & count <= _T_27 ? _GEN_154 : L0Memory_25; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_255 = count >= 10'h1 & count <= _T_27 ? _GEN_155 : L0Memory_26; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_256 = count >= 10'h1 & count <= _T_27 ? _GEN_156 : L0Memory_27; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_257 = count >= 10'h1 & count <= _T_27 ? _GEN_157 : L0Memory_28; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_258 = count >= 10'h1 & count <= _T_27 ? _GEN_158 : L0Memory_29; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_259 = count >= 10'h1 & count <= _T_27 ? _GEN_159 : L0Memory_30; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_260 = count >= 10'h1 & count <= _T_27 ? _GEN_160 : L0Memory_31; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_261 = count >= 10'h1 & count <= _T_27 ? _GEN_161 : L0Memory_32; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_262 = count >= 10'h1 & count <= _T_27 ? _GEN_162 : L0Memory_33; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_263 = count >= 10'h1 & count <= _T_27 ? _GEN_163 : L0Memory_34; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_264 = count >= 10'h1 & count <= _T_27 ? _GEN_164 : L0Memory_35; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_265 = count >= 10'h1 & count <= _T_27 ? _GEN_165 : L0Memory_36; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_266 = count >= 10'h1 & count <= _T_27 ? _GEN_166 : L0Memory_37; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_267 = count >= 10'h1 & count <= _T_27 ? _GEN_167 : L0Memory_38; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_268 = count >= 10'h1 & count <= _T_27 ? _GEN_168 : L0Memory_39; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_269 = count >= 10'h1 & count <= _T_27 ? _GEN_169 : L0Memory_40; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_270 = count >= 10'h1 & count <= _T_27 ? _GEN_170 : L0Memory_41; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_271 = count >= 10'h1 & count <= _T_27 ? _GEN_171 : L0Memory_42; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_272 = count >= 10'h1 & count <= _T_27 ? _GEN_172 : L0Memory_43; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_273 = count >= 10'h1 & count <= _T_27 ? _GEN_173 : L0Memory_44; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_274 = count >= 10'h1 & count <= _T_27 ? _GEN_174 : L0Memory_45; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_275 = count >= 10'h1 & count <= _T_27 ? _GEN_175 : L0Memory_46; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_276 = count >= 10'h1 & count <= _T_27 ? _GEN_176 : L0Memory_47; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_277 = count >= 10'h1 & count <= _T_27 ? _GEN_177 : L0Memory_48; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_278 = count >= 10'h1 & count <= _T_27 ? _GEN_178 : L0Memory_49; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_279 = count >= 10'h1 & count <= _T_27 ? _GEN_179 : L0Memory_50; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_280 = count >= 10'h1 & count <= _T_27 ? _GEN_180 : L0Memory_51; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_281 = count >= 10'h1 & count <= _T_27 ? _GEN_181 : L0Memory_52; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_282 = count >= 10'h1 & count <= _T_27 ? _GEN_182 : L0Memory_53; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_283 = count >= 10'h1 & count <= _T_27 ? _GEN_183 : L0Memory_54; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_284 = count >= 10'h1 & count <= _T_27 ? _GEN_184 : L0Memory_55; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_285 = count >= 10'h1 & count <= _T_27 ? _GEN_185 : L0Memory_56; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_286 = count >= 10'h1 & count <= _T_27 ? _GEN_186 : L0Memory_57; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_287 = count >= 10'h1 & count <= _T_27 ? _GEN_187 : L0Memory_58; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_288 = count >= 10'h1 & count <= _T_27 ? _GEN_188 : L0Memory_59; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_289 = count >= 10'h1 & count <= _T_27 ? _GEN_189 : L0Memory_60; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_290 = count >= 10'h1 & count <= _T_27 ? _GEN_190 : L0Memory_61; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_291 = count >= 10'h1 & count <= _T_27 ? _GEN_191 : L0Memory_62; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_292 = count >= 10'h1 & count <= _T_27 ? _GEN_192 : L0Memory_63; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_293 = count >= 10'h1 & count <= _T_27 ? _GEN_193 : L0Memory_64; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_294 = count >= 10'h1 & count <= _T_27 ? _GEN_194 : L0Memory_65; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_295 = count >= 10'h1 & count <= _T_27 ? _GEN_195 : L0Memory_66; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_296 = count >= 10'h1 & count <= _T_27 ? _GEN_196 : L0Memory_67; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_297 = count >= 10'h1 & count <= _T_27 ? _GEN_197 : L0Memory_68; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_298 = count >= 10'h1 & count <= _T_27 ? _GEN_198 : L0Memory_69; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_299 = count >= 10'h1 & count <= _T_27 ? _GEN_199 : L0Memory_70; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_300 = count >= 10'h1 & count <= _T_27 ? _GEN_200 : L0Memory_71; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_301 = count >= 10'h1 & count <= _T_27 ? _GEN_201 : L0Memory_72; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_302 = count >= 10'h1 & count <= _T_27 ? _GEN_202 : L0Memory_73; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_303 = count >= 10'h1 & count <= _T_27 ? _GEN_203 : L0Memory_74; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_304 = count >= 10'h1 & count <= _T_27 ? _GEN_204 : L0Memory_75; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_305 = count >= 10'h1 & count <= _T_27 ? _GEN_205 : L0Memory_76; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_306 = count >= 10'h1 & count <= _T_27 ? _GEN_206 : L0Memory_77; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_307 = count >= 10'h1 & count <= _T_27 ? _GEN_207 : L0Memory_78; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_308 = count >= 10'h1 & count <= _T_27 ? _GEN_208 : L0Memory_79; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_309 = count >= 10'h1 & count <= _T_27 ? _GEN_209 : L0Memory_80; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_310 = count >= 10'h1 & count <= _T_27 ? _GEN_210 : L0Memory_81; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_311 = count >= 10'h1 & count <= _T_27 ? _GEN_211 : L0Memory_82; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_312 = count >= 10'h1 & count <= _T_27 ? _GEN_212 : L0Memory_83; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_313 = count >= 10'h1 & count <= _T_27 ? _GEN_213 : L0Memory_84; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_314 = count >= 10'h1 & count <= _T_27 ? _GEN_214 : L0Memory_85; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_315 = count >= 10'h1 & count <= _T_27 ? _GEN_215 : L0Memory_86; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_316 = count >= 10'h1 & count <= _T_27 ? _GEN_216 : L0Memory_87; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_317 = count >= 10'h1 & count <= _T_27 ? _GEN_217 : L0Memory_88; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_318 = count >= 10'h1 & count <= _T_27 ? _GEN_218 : L0Memory_89; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_319 = count >= 10'h1 & count <= _T_27 ? _GEN_219 : L0Memory_90; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_320 = count >= 10'h1 & count <= _T_27 ? _GEN_220 : L0Memory_91; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_321 = count >= 10'h1 & count <= _T_27 ? _GEN_221 : L0Memory_92; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_322 = count >= 10'h1 & count <= _T_27 ? _GEN_222 : L0Memory_93; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_323 = count >= 10'h1 & count <= _T_27 ? _GEN_223 : L0Memory_94; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_324 = count >= 10'h1 & count <= _T_27 ? _GEN_224 : L0Memory_95; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_325 = count >= 10'h1 & count <= _T_27 ? _GEN_225 : L0Memory_96; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_326 = count >= 10'h1 & count <= _T_27 ? _GEN_226 : L0Memory_97; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_327 = count >= 10'h1 & count <= _T_27 ? _GEN_227 : L0Memory_98; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_328 = count >= 10'h1 & count <= _T_27 ? _GEN_228 : L0Memory_99; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [5:0] _GEN_329 = count >= 10'h1 & count <= _T_27 ? _L0Index_T_2 : _GEN_128; // @[PEArray.scala 198:59 PEArray.scala 200:17]
  wire [9:0] _GEN_330 = count == count_max ? 10'h0 : _GEN_127; // @[PEArray.scala 202:32 PEArray.scala 203:15]
  wire [2:0] _GEN_331 = count == count_max ? 3'h0 : state; // @[PEArray.scala 202:32 PEArray.scala 204:15 PEArray.scala 100:22]
  wire [9:0] _GEN_865 = {{4'd0}, GRU_out_width}; // @[PEArray.scala 220:19]
  wire [9:0] _GEN_0 = count % _GEN_865; // @[PEArray.scala 220:19]
  wire [5:0] _T_36 = _GEN_0[5:0]; // @[PEArray.scala 220:19]
  wire [5:0] _T_38 = GRU_out_width - 6'h1; // @[PEArray.scala 220:55]
  wire [5:0] _GEN_334 = _T_36 == _T_38 ? _L0Index_T_2 : L0index_begin; // @[PEArray.scala 220:62 PEArray.scala 221:17 PEArray.scala 214:15]
  wire [5:0] _GEN_346 = _T_41 ? _GEN_334 : L0Index; // @[Conditional.scala 39:67 PEArray.scala 39:24]
  wire [9:0] _GEN_347 = _T_41 ? _GEN_330 : count; // @[Conditional.scala 39:67 PEArray.scala 101:22]
  wire [2:0] _GEN_348 = _T_41 ? _GEN_331 : state; // @[Conditional.scala 39:67 PEArray.scala 100:22]
  wire [5:0] _GEN_353 = _T_31 ? _GEN_334 : _GEN_346; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_354 = _T_31 ? _GEN_330 : _GEN_347; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_355 = _T_31 ? _GEN_331 : _GEN_348; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_356 = _T_22 ? _GEN_330 : _GEN_354; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_357 = _T_22 ? _GEN_329 : _GEN_353; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_458 = _T_22 ? _GEN_331 : _GEN_355; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_690 = _T_3 ? _GEN_118 : {{2'd0}, GRU_out_width}; // @[Conditional.scala 40:58 PEArray.scala 104:26]
  FP16MulAdder FP16MAC ( // @[PEArray.scala 72:23]
    .io_a(FP16MAC_io_a),
    .io_b(FP16MAC_io_b),
    .io_c(FP16MAC_io_c),
    .io_out(FP16MAC_io_out)
  );
  assign io_ToRightPE = mux3out_reg; // @[PEArray.scala 95:16]
  assign io_ToBelowPE = mux2out_reg; // @[PEArray.scala 94:16]
  assign FP16MAC_io_a = sel1 ? io_FromL1 : io_FromLeftPE; // @[PEArray.scala 50:14 PEArray.scala 50:23 PEArray.scala 51:24]
  assign FP16MAC_io_b = sel5 ? mux4out : _GEN_105; // @[PEArray.scala 77:13 PEArray.scala 78:18 PEArray.scala 81:18]
  assign FP16MAC_io_c = sel5 ? _GEN_105 : mux4out; // @[PEArray.scala 77:13 PEArray.scala 79:18 PEArray.scala 82:18]
  always @(posedge clock) begin
    if (reset) begin // @[PEArray.scala 39:24]
      L0Index <= 6'h0; // @[PEArray.scala 39:24]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h2; // @[PEArray.scala 159:15]
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h6; // @[PEArray.scala 181:15]
      end else begin
        L0Index <= _GEN_357;
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_0 <= _GEN_229;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_1 <= _GEN_230;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_2 <= _GEN_231;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_3 <= _GEN_232;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_4 <= _GEN_233;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_5 <= _GEN_234;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_6 <= _GEN_235;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_7 <= _GEN_236;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_8 <= _GEN_237;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_9 <= _GEN_238;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_10 <= _GEN_239;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_11 <= _GEN_240;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_12 <= _GEN_241;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_13 <= _GEN_242;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_14 <= _GEN_243;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_15 <= _GEN_244;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_16 <= _GEN_245;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_17 <= _GEN_246;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_18 <= _GEN_247;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_19 <= _GEN_248;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_20 <= _GEN_249;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_21 <= _GEN_250;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_22 <= _GEN_251;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_23 <= _GEN_252;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_24 <= _GEN_253;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_25 <= _GEN_254;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_26 <= _GEN_255;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_27 <= _GEN_256;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_28 <= _GEN_257;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_29 <= _GEN_258;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_30 <= _GEN_259;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_31 <= _GEN_260;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_32 <= _GEN_261;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_33 <= _GEN_262;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_34 <= _GEN_263;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_35 <= _GEN_264;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_36 <= _GEN_265;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_37 <= _GEN_266;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_38 <= _GEN_267;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_39 <= _GEN_268;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_40 <= _GEN_269;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_41 <= _GEN_270;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_42 <= _GEN_271;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_43 <= _GEN_272;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_44 <= _GEN_273;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_45 <= _GEN_274;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_46 <= _GEN_275;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_47 <= _GEN_276;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_48 <= _GEN_277;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_49 <= _GEN_278;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_50 <= _GEN_279;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_51 <= _GEN_280;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_52 <= _GEN_281;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_53 <= _GEN_282;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_54 <= _GEN_283;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_55 <= _GEN_284;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_56 <= _GEN_285;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_57 <= _GEN_286;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_58 <= _GEN_287;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_59 <= _GEN_288;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_60 <= _GEN_289;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_61 <= _GEN_290;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_62 <= _GEN_291;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_63 <= _GEN_292;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_64 <= _GEN_293;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_65 <= _GEN_294;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_66 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_67 <= _GEN_296;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_68 <= _GEN_297;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_69 <= _GEN_298;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_70 <= _GEN_299;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_71 <= _GEN_300;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_72 <= _GEN_301;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_73 <= _GEN_302;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_74 <= _GEN_303;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_75 <= _GEN_304;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_76 <= _GEN_305;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_77 <= _GEN_306;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_78 <= _GEN_307;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_79 <= _GEN_308;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_80 <= _GEN_309;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_81 <= _GEN_310;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_82 <= _GEN_311;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_83 <= _GEN_312;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_84 <= _GEN_313;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_85 <= _GEN_314;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_86 <= _GEN_315;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_87 <= _GEN_316;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_88 <= _GEN_317;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_89 <= _GEN_318;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_90 <= _GEN_319;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_91 <= _GEN_320;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_92 <= _GEN_321;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_93 <= _GEN_322;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_94 <= _GEN_323;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_95 <= _GEN_324;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_96 <= _GEN_325;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_97 <= _GEN_326;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_98 <= _GEN_327;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_99 <= _GEN_328;
          end
        end
      end
    end
    if (reset) begin // @[PEArray.scala 100:22]
      state <= 3'h0; // @[PEArray.scala 100:22]
    end else if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[8]) begin // @[PEArray.scala 116:57]
        if (_T_6) begin // @[Conditional.scala 40:58]
          state <= 3'h0; // @[PEArray.scala 120:19]
        end else begin
          state <= _GEN_113;
        end
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      if (count == 10'h33) begin // @[PEArray.scala 164:27]
        state <= 3'h0; // @[PEArray.scala 166:15]
      end
    end else if (_T_16) begin // @[Conditional.scala 39:67]
      state <= _GEN_126;
    end else begin
      state <= _GEN_458;
    end
    if (reset) begin // @[PEArray.scala 90:28]
      mux2out_reg <= 16'h0; // @[PEArray.scala 90:28]
    end else begin
      mux2out_reg <= MAC_out; // @[PEArray.scala 90:28]
    end
    if (reset) begin // @[PEArray.scala 91:28]
      mux3out_reg <= 16'h0; // @[PEArray.scala 91:28]
    end else if (sel3) begin // @[PEArray.scala 56:14]
      mux3out_reg <= MAC_out; // @[PEArray.scala 56:23]
    end else if (sel1) begin // @[PEArray.scala 50:14]
      mux3out_reg <= io_FromL1; // @[PEArray.scala 50:23]
    end else begin
      mux3out_reg <= io_FromLeftPE; // @[PEArray.scala 51:24]
    end
    if (reset) begin // @[PEArray.scala 101:22]
      count <= 10'h0; // @[PEArray.scala 101:22]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        if (count == 10'h33) begin // @[PEArray.scala 164:27]
          count <= 10'h0; // @[PEArray.scala 165:15]
        end else begin
          count <= _GEN_120;
        end
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        count <= _GEN_125;
      end else begin
        count <= _GEN_356;
      end
    end
    if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[8]) begin // @[PEArray.scala 116:57]
        count_max <= io_control_signal_count; // @[PEArray.scala 143:19]
      end
    end
    if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[8]) begin // @[PEArray.scala 116:57]
        L0index_begin <= io_control_signal_L0index; // @[PEArray.scala 144:23]
      end
    end
    GRU_out_width <= _GEN_690[5:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  L0Index = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  L0Memory_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  L0Memory_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  L0Memory_2 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  L0Memory_3 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  L0Memory_4 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  L0Memory_5 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  L0Memory_6 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  L0Memory_7 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  L0Memory_8 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  L0Memory_9 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  L0Memory_10 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  L0Memory_11 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  L0Memory_12 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  L0Memory_13 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  L0Memory_14 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  L0Memory_15 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  L0Memory_16 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  L0Memory_17 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  L0Memory_18 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  L0Memory_19 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  L0Memory_20 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  L0Memory_21 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  L0Memory_22 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  L0Memory_23 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  L0Memory_24 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  L0Memory_25 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  L0Memory_26 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  L0Memory_27 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  L0Memory_28 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  L0Memory_29 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  L0Memory_30 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  L0Memory_31 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  L0Memory_32 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  L0Memory_33 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  L0Memory_34 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  L0Memory_35 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  L0Memory_36 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  L0Memory_37 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  L0Memory_38 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  L0Memory_39 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  L0Memory_40 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  L0Memory_41 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  L0Memory_42 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  L0Memory_43 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  L0Memory_44 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  L0Memory_45 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  L0Memory_46 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  L0Memory_47 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  L0Memory_48 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  L0Memory_49 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  L0Memory_50 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  L0Memory_51 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  L0Memory_52 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  L0Memory_53 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  L0Memory_54 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  L0Memory_55 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  L0Memory_56 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  L0Memory_57 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  L0Memory_58 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  L0Memory_59 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  L0Memory_60 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  L0Memory_61 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  L0Memory_62 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  L0Memory_63 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  L0Memory_64 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  L0Memory_65 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  L0Memory_66 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  L0Memory_67 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  L0Memory_68 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  L0Memory_69 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  L0Memory_70 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  L0Memory_71 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  L0Memory_72 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  L0Memory_73 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  L0Memory_74 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  L0Memory_75 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  L0Memory_76 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  L0Memory_77 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  L0Memory_78 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  L0Memory_79 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  L0Memory_80 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  L0Memory_81 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  L0Memory_82 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  L0Memory_83 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  L0Memory_84 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  L0Memory_85 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  L0Memory_86 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  L0Memory_87 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  L0Memory_88 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  L0Memory_89 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  L0Memory_90 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  L0Memory_91 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  L0Memory_92 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  L0Memory_93 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  L0Memory_94 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  L0Memory_95 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  L0Memory_96 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  L0Memory_97 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  L0Memory_98 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  L0Memory_99 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  state = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  mux2out_reg = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  mux3out_reg = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  count = _RAND_104[9:0];
  _RAND_105 = {1{`RANDOM}};
  count_max = _RAND_105[9:0];
  _RAND_106 = {1{`RANDOM}};
  L0index_begin = _RAND_106[5:0];
  _RAND_107 = {1{`RANDOM}};
  GRU_out_width = _RAND_107[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PE_12(
  input         clock,
  input         reset,
  input  [15:0] io_FromAbovePE,
  input  [15:0] io_FromLeftPE,
  input  [15:0] io_FromL1,
  input  [11:0] io_control_signal_mask,
  output [15:0] io_ToRightPE,
  output [15:0] io_ToBelowPE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] FP16MAC_io_a; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_b; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_c; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_out; // @[PEArray.scala 72:23]
  reg [5:0] L0Index; // @[PEArray.scala 39:24]
  reg [15:0] L0Memory_0; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_1; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_2; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_3; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_4; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_5; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_6; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_7; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_8; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_9; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_10; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_11; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_12; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_13; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_14; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_15; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_16; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_17; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_18; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_19; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_20; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_21; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_22; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_23; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_24; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_25; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_26; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_27; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_28; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_29; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_30; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_31; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_32; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_33; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_34; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_35; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_36; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_37; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_38; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_39; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_40; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_41; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_42; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_43; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_44; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_45; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_46; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_47; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_48; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_49; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_50; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_51; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_52; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_53; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_54; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_55; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_56; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_57; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_58; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_59; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_60; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_61; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_62; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_63; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_64; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_65; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_66; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_67; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_68; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_69; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_70; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_71; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_72; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_73; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_74; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_75; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_76; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_77; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_78; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_79; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_80; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_81; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_82; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_83; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_84; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_85; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_86; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_87; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_88; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_89; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_90; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_91; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_92; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_93; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_94; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_95; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_96; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_97; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_98; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_99; // @[PEArray.scala 40:21]
  reg [2:0] state; // @[PEArray.scala 100:22]
  wire  _T_3 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_12 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_16 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_22 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_31 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_41 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_342 = _T_41 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 231:12 PEArray.scala 32:8]
  wire  _GEN_349 = _T_31 ? 1'h0 : _GEN_342; // @[Conditional.scala 39:67 PEArray.scala 208:12]
  wire  _GEN_459 = _T_22 | _GEN_349; // @[Conditional.scala 39:67 PEArray.scala 32:8]
  wire  _GEN_463 = _T_16 ? 1'h0 : _GEN_459; // @[Conditional.scala 39:67]
  wire  _GEN_572 = _T_12 | _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 149:12]
  wire  sel1 = _T_3 | _GEN_572; // @[Conditional.scala 40:58 PEArray.scala 108:12]
  wire [15:0] MAC_out = FP16MAC_io_out; // @[PEArray.scala 47:21 PEArray.scala 85:11]
  wire  _GEN_465 = _T_16 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 177:12]
  wire  _GEN_580 = _T_12 | _GEN_465; // @[Conditional.scala 39:67 PEArray.scala 34:8]
  wire  sel3 = _T_3 | _GEN_580; // @[Conditional.scala 40:58 PEArray.scala 110:12]
  wire [1:0] _GEN_344 = _T_41 ? 2'h2 : 2'h0; // @[Conditional.scala 39:67 PEArray.scala 233:12 PEArray.scala 35:8]
  wire [1:0] _GEN_351 = _T_31 ? 2'h2 : _GEN_344; // @[Conditional.scala 39:67 PEArray.scala 210:12]
  wire [1:0] _GEN_461 = _T_22 ? 2'h0 : _GEN_351; // @[Conditional.scala 39:67 PEArray.scala 35:8]
  wire [1:0] _GEN_466 = _T_16 ? 2'h0 : _GEN_461; // @[Conditional.scala 39:67 PEArray.scala 178:12]
  wire [1:0] _GEN_574 = _T_12 ? 2'h0 : _GEN_466; // @[Conditional.scala 39:67]
  wire [1:0] sel4 = _T_3 ? 2'h0 : _GEN_574; // @[Conditional.scala 40:58 PEArray.scala 111:12]
  wire [15:0] _GEN_3 = sel4 == 2'h2 ? io_FromL1 : 16'h0; // @[PEArray.scala 65:28 PEArray.scala 66:15 PEArray.scala 69:15]
  wire [15:0] _GEN_4 = sel4 == 2'h1 ? io_FromAbovePE : _GEN_3; // @[PEArray.scala 62:28 PEArray.scala 63:15]
  wire [15:0] mux4out = sel4 == 2'h0 ? 16'h0 : _GEN_4; // @[PEArray.scala 59:22 PEArray.scala 60:13]
  wire [15:0] _GEN_7 = 6'h1 == L0Index ? L0Memory_1 : L0Memory_0; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_8 = 6'h2 == L0Index ? L0Memory_2 : _GEN_7; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_9 = 6'h3 == L0Index ? L0Memory_3 : _GEN_8; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_10 = 6'h4 == L0Index ? L0Memory_4 : _GEN_9; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_11 = 6'h5 == L0Index ? L0Memory_5 : _GEN_10; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_12 = 6'h6 == L0Index ? L0Memory_6 : _GEN_11; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_13 = 6'h7 == L0Index ? L0Memory_7 : _GEN_12; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_14 = 6'h8 == L0Index ? L0Memory_8 : _GEN_13; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_15 = 6'h9 == L0Index ? L0Memory_9 : _GEN_14; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_16 = 6'ha == L0Index ? L0Memory_10 : _GEN_15; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_17 = 6'hb == L0Index ? L0Memory_11 : _GEN_16; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_18 = 6'hc == L0Index ? L0Memory_12 : _GEN_17; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_19 = 6'hd == L0Index ? L0Memory_13 : _GEN_18; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_20 = 6'he == L0Index ? L0Memory_14 : _GEN_19; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_21 = 6'hf == L0Index ? L0Memory_15 : _GEN_20; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_22 = 6'h10 == L0Index ? L0Memory_16 : _GEN_21; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_23 = 6'h11 == L0Index ? L0Memory_17 : _GEN_22; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_24 = 6'h12 == L0Index ? L0Memory_18 : _GEN_23; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_25 = 6'h13 == L0Index ? L0Memory_19 : _GEN_24; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_26 = 6'h14 == L0Index ? L0Memory_20 : _GEN_25; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_27 = 6'h15 == L0Index ? L0Memory_21 : _GEN_26; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_28 = 6'h16 == L0Index ? L0Memory_22 : _GEN_27; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_29 = 6'h17 == L0Index ? L0Memory_23 : _GEN_28; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_30 = 6'h18 == L0Index ? L0Memory_24 : _GEN_29; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_31 = 6'h19 == L0Index ? L0Memory_25 : _GEN_30; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_32 = 6'h1a == L0Index ? L0Memory_26 : _GEN_31; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_33 = 6'h1b == L0Index ? L0Memory_27 : _GEN_32; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_34 = 6'h1c == L0Index ? L0Memory_28 : _GEN_33; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_35 = 6'h1d == L0Index ? L0Memory_29 : _GEN_34; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_36 = 6'h1e == L0Index ? L0Memory_30 : _GEN_35; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_37 = 6'h1f == L0Index ? L0Memory_31 : _GEN_36; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_38 = 6'h20 == L0Index ? L0Memory_32 : _GEN_37; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_39 = 6'h21 == L0Index ? L0Memory_33 : _GEN_38; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_40 = 6'h22 == L0Index ? L0Memory_34 : _GEN_39; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_41 = 6'h23 == L0Index ? L0Memory_35 : _GEN_40; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_42 = 6'h24 == L0Index ? L0Memory_36 : _GEN_41; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_43 = 6'h25 == L0Index ? L0Memory_37 : _GEN_42; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_44 = 6'h26 == L0Index ? L0Memory_38 : _GEN_43; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_45 = 6'h27 == L0Index ? L0Memory_39 : _GEN_44; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_46 = 6'h28 == L0Index ? L0Memory_40 : _GEN_45; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_47 = 6'h29 == L0Index ? L0Memory_41 : _GEN_46; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_48 = 6'h2a == L0Index ? L0Memory_42 : _GEN_47; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_49 = 6'h2b == L0Index ? L0Memory_43 : _GEN_48; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_50 = 6'h2c == L0Index ? L0Memory_44 : _GEN_49; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_51 = 6'h2d == L0Index ? L0Memory_45 : _GEN_50; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_52 = 6'h2e == L0Index ? L0Memory_46 : _GEN_51; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_53 = 6'h2f == L0Index ? L0Memory_47 : _GEN_52; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_54 = 6'h30 == L0Index ? L0Memory_48 : _GEN_53; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_55 = 6'h31 == L0Index ? L0Memory_49 : _GEN_54; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_56 = 6'h32 == L0Index ? L0Memory_50 : _GEN_55; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_57 = 6'h33 == L0Index ? L0Memory_51 : _GEN_56; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_58 = 6'h34 == L0Index ? L0Memory_52 : _GEN_57; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_59 = 6'h35 == L0Index ? L0Memory_53 : _GEN_58; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_60 = 6'h36 == L0Index ? L0Memory_54 : _GEN_59; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_61 = 6'h37 == L0Index ? L0Memory_55 : _GEN_60; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_62 = 6'h38 == L0Index ? L0Memory_56 : _GEN_61; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_63 = 6'h39 == L0Index ? L0Memory_57 : _GEN_62; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_64 = 6'h3a == L0Index ? L0Memory_58 : _GEN_63; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_65 = 6'h3b == L0Index ? L0Memory_59 : _GEN_64; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_66 = 6'h3c == L0Index ? L0Memory_60 : _GEN_65; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_67 = 6'h3d == L0Index ? L0Memory_61 : _GEN_66; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_68 = 6'h3e == L0Index ? L0Memory_62 : _GEN_67; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_69 = 6'h3f == L0Index ? L0Memory_63 : _GEN_68; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [6:0] _GEN_793 = {{1'd0}, L0Index}; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_70 = 7'h40 == _GEN_793 ? L0Memory_64 : _GEN_69; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_71 = 7'h41 == _GEN_793 ? L0Memory_65 : _GEN_70; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_72 = 7'h42 == _GEN_793 ? L0Memory_66 : _GEN_71; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_73 = 7'h43 == _GEN_793 ? L0Memory_67 : _GEN_72; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_74 = 7'h44 == _GEN_793 ? L0Memory_68 : _GEN_73; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_75 = 7'h45 == _GEN_793 ? L0Memory_69 : _GEN_74; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_76 = 7'h46 == _GEN_793 ? L0Memory_70 : _GEN_75; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_77 = 7'h47 == _GEN_793 ? L0Memory_71 : _GEN_76; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_78 = 7'h48 == _GEN_793 ? L0Memory_72 : _GEN_77; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_79 = 7'h49 == _GEN_793 ? L0Memory_73 : _GEN_78; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_80 = 7'h4a == _GEN_793 ? L0Memory_74 : _GEN_79; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_81 = 7'h4b == _GEN_793 ? L0Memory_75 : _GEN_80; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_82 = 7'h4c == _GEN_793 ? L0Memory_76 : _GEN_81; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_83 = 7'h4d == _GEN_793 ? L0Memory_77 : _GEN_82; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_84 = 7'h4e == _GEN_793 ? L0Memory_78 : _GEN_83; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_85 = 7'h4f == _GEN_793 ? L0Memory_79 : _GEN_84; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_86 = 7'h50 == _GEN_793 ? L0Memory_80 : _GEN_85; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_87 = 7'h51 == _GEN_793 ? L0Memory_81 : _GEN_86; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_88 = 7'h52 == _GEN_793 ? L0Memory_82 : _GEN_87; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_89 = 7'h53 == _GEN_793 ? L0Memory_83 : _GEN_88; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_90 = 7'h54 == _GEN_793 ? L0Memory_84 : _GEN_89; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_91 = 7'h55 == _GEN_793 ? L0Memory_85 : _GEN_90; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_92 = 7'h56 == _GEN_793 ? L0Memory_86 : _GEN_91; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_93 = 7'h57 == _GEN_793 ? L0Memory_87 : _GEN_92; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_94 = 7'h58 == _GEN_793 ? L0Memory_88 : _GEN_93; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_95 = 7'h59 == _GEN_793 ? L0Memory_89 : _GEN_94; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_96 = 7'h5a == _GEN_793 ? L0Memory_90 : _GEN_95; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_97 = 7'h5b == _GEN_793 ? L0Memory_91 : _GEN_96; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_98 = 7'h5c == _GEN_793 ? L0Memory_92 : _GEN_97; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_99 = 7'h5d == _GEN_793 ? L0Memory_93 : _GEN_98; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_100 = 7'h5e == _GEN_793 ? L0Memory_94 : _GEN_99; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_101 = 7'h5f == _GEN_793 ? L0Memory_95 : _GEN_100; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_102 = 7'h60 == _GEN_793 ? L0Memory_96 : _GEN_101; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_103 = 7'h61 == _GEN_793 ? L0Memory_97 : _GEN_102; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_104 = 7'h62 == _GEN_793 ? L0Memory_98 : _GEN_103; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_105 = 7'h63 == _GEN_793 ? L0Memory_99 : _GEN_104; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire  _GEN_575 = _T_12 ? 1'h0 : _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 157:12]
  wire  sel5 = _T_3 ? 1'h0 : _GEN_575; // @[Conditional.scala 40:58 PEArray.scala 112:12]
  reg [15:0] mux2out_reg; // @[PEArray.scala 90:28]
  reg [15:0] mux3out_reg; // @[PEArray.scala 91:28]
  reg [9:0] count; // @[PEArray.scala 101:22]
  reg [5:0] GRU_out_width; // @[PEArray.scala 104:26]
  wire [7:0] _GEN_118 = io_control_signal_mask[7] ? 8'h0 : {{2'd0}, GRU_out_width}; // @[PEArray.scala 116:57 PEArray.scala 145:23 PEArray.scala 104:26]
  wire [9:0] _count_T_1 = count + 10'h1; // @[PEArray.scala 162:24]
  wire [9:0] _GEN_120 = count != 10'h33 ? _count_T_1 : count; // @[PEArray.scala 161:27 PEArray.scala 162:15 PEArray.scala 101:22]
  wire [9:0] _GEN_124 = count != 10'h188 ? _count_T_1 : count; // @[PEArray.scala 183:28 PEArray.scala 184:15 PEArray.scala 101:22]
  wire [9:0] _GEN_125 = count == 10'h188 ? 10'h0 : _GEN_124; // @[PEArray.scala 186:28 PEArray.scala 187:15]
  wire [2:0] _GEN_126 = count == 10'h188 ? 3'h0 : state; // @[PEArray.scala 186:28 PEArray.scala 188:15 PEArray.scala 100:22]
  wire [9:0] _GEN_127 = count != 10'h0 ? _count_T_1 : count; // @[PEArray.scala 192:32 PEArray.scala 193:15 PEArray.scala 101:22]
  wire  _T_24 = count == 10'h0; // @[PEArray.scala 195:18]
  wire [5:0] _GEN_128 = count == 10'h0 ? 6'h0 : L0Index; // @[PEArray.scala 195:26 PEArray.scala 196:17 PEArray.scala 39:24]
  wire [9:0] _T_27 = 10'h0 - 10'h1; // @[PEArray.scala 198:51]
  wire [15:0] _GEN_129 = 6'h0 == L0Index ? io_FromL1 : L0Memory_0; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_130 = 6'h1 == L0Index ? io_FromL1 : L0Memory_1; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_131 = 6'h2 == L0Index ? io_FromL1 : L0Memory_2; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_132 = 6'h3 == L0Index ? io_FromL1 : L0Memory_3; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_133 = 6'h4 == L0Index ? io_FromL1 : L0Memory_4; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_134 = 6'h5 == L0Index ? io_FromL1 : L0Memory_5; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_135 = 6'h6 == L0Index ? io_FromL1 : L0Memory_6; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_136 = 6'h7 == L0Index ? io_FromL1 : L0Memory_7; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_137 = 6'h8 == L0Index ? io_FromL1 : L0Memory_8; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_138 = 6'h9 == L0Index ? io_FromL1 : L0Memory_9; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_139 = 6'ha == L0Index ? io_FromL1 : L0Memory_10; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_140 = 6'hb == L0Index ? io_FromL1 : L0Memory_11; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_141 = 6'hc == L0Index ? io_FromL1 : L0Memory_12; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_142 = 6'hd == L0Index ? io_FromL1 : L0Memory_13; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_143 = 6'he == L0Index ? io_FromL1 : L0Memory_14; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_144 = 6'hf == L0Index ? io_FromL1 : L0Memory_15; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_145 = 6'h10 == L0Index ? io_FromL1 : L0Memory_16; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_146 = 6'h11 == L0Index ? io_FromL1 : L0Memory_17; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_147 = 6'h12 == L0Index ? io_FromL1 : L0Memory_18; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_148 = 6'h13 == L0Index ? io_FromL1 : L0Memory_19; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_149 = 6'h14 == L0Index ? io_FromL1 : L0Memory_20; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_150 = 6'h15 == L0Index ? io_FromL1 : L0Memory_21; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_151 = 6'h16 == L0Index ? io_FromL1 : L0Memory_22; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_152 = 6'h17 == L0Index ? io_FromL1 : L0Memory_23; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_153 = 6'h18 == L0Index ? io_FromL1 : L0Memory_24; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_154 = 6'h19 == L0Index ? io_FromL1 : L0Memory_25; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_155 = 6'h1a == L0Index ? io_FromL1 : L0Memory_26; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_156 = 6'h1b == L0Index ? io_FromL1 : L0Memory_27; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_157 = 6'h1c == L0Index ? io_FromL1 : L0Memory_28; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_158 = 6'h1d == L0Index ? io_FromL1 : L0Memory_29; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_159 = 6'h1e == L0Index ? io_FromL1 : L0Memory_30; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_160 = 6'h1f == L0Index ? io_FromL1 : L0Memory_31; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_161 = 6'h20 == L0Index ? io_FromL1 : L0Memory_32; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_162 = 6'h21 == L0Index ? io_FromL1 : L0Memory_33; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_163 = 6'h22 == L0Index ? io_FromL1 : L0Memory_34; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_164 = 6'h23 == L0Index ? io_FromL1 : L0Memory_35; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_165 = 6'h24 == L0Index ? io_FromL1 : L0Memory_36; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_166 = 6'h25 == L0Index ? io_FromL1 : L0Memory_37; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_167 = 6'h26 == L0Index ? io_FromL1 : L0Memory_38; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_168 = 6'h27 == L0Index ? io_FromL1 : L0Memory_39; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_169 = 6'h28 == L0Index ? io_FromL1 : L0Memory_40; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_170 = 6'h29 == L0Index ? io_FromL1 : L0Memory_41; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_171 = 6'h2a == L0Index ? io_FromL1 : L0Memory_42; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_172 = 6'h2b == L0Index ? io_FromL1 : L0Memory_43; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_173 = 6'h2c == L0Index ? io_FromL1 : L0Memory_44; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_174 = 6'h2d == L0Index ? io_FromL1 : L0Memory_45; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_175 = 6'h2e == L0Index ? io_FromL1 : L0Memory_46; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_176 = 6'h2f == L0Index ? io_FromL1 : L0Memory_47; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_177 = 6'h30 == L0Index ? io_FromL1 : L0Memory_48; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_178 = 6'h31 == L0Index ? io_FromL1 : L0Memory_49; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_179 = 6'h32 == L0Index ? io_FromL1 : L0Memory_50; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_180 = 6'h33 == L0Index ? io_FromL1 : L0Memory_51; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_181 = 6'h34 == L0Index ? io_FromL1 : L0Memory_52; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_182 = 6'h35 == L0Index ? io_FromL1 : L0Memory_53; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_183 = 6'h36 == L0Index ? io_FromL1 : L0Memory_54; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_184 = 6'h37 == L0Index ? io_FromL1 : L0Memory_55; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_185 = 6'h38 == L0Index ? io_FromL1 : L0Memory_56; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_186 = 6'h39 == L0Index ? io_FromL1 : L0Memory_57; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_187 = 6'h3a == L0Index ? io_FromL1 : L0Memory_58; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_188 = 6'h3b == L0Index ? io_FromL1 : L0Memory_59; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_189 = 6'h3c == L0Index ? io_FromL1 : L0Memory_60; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_190 = 6'h3d == L0Index ? io_FromL1 : L0Memory_61; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_191 = 6'h3e == L0Index ? io_FromL1 : L0Memory_62; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_192 = 6'h3f == L0Index ? io_FromL1 : L0Memory_63; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_193 = 7'h40 == _GEN_793 ? io_FromL1 : L0Memory_64; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_194 = 7'h41 == _GEN_793 ? io_FromL1 : L0Memory_65; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_195 = 7'h42 == _GEN_793 ? io_FromL1 : L0Memory_66; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_196 = 7'h43 == _GEN_793 ? io_FromL1 : L0Memory_67; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_197 = 7'h44 == _GEN_793 ? io_FromL1 : L0Memory_68; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_198 = 7'h45 == _GEN_793 ? io_FromL1 : L0Memory_69; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_199 = 7'h46 == _GEN_793 ? io_FromL1 : L0Memory_70; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_200 = 7'h47 == _GEN_793 ? io_FromL1 : L0Memory_71; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_201 = 7'h48 == _GEN_793 ? io_FromL1 : L0Memory_72; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_202 = 7'h49 == _GEN_793 ? io_FromL1 : L0Memory_73; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_203 = 7'h4a == _GEN_793 ? io_FromL1 : L0Memory_74; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_204 = 7'h4b == _GEN_793 ? io_FromL1 : L0Memory_75; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_205 = 7'h4c == _GEN_793 ? io_FromL1 : L0Memory_76; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_206 = 7'h4d == _GEN_793 ? io_FromL1 : L0Memory_77; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_207 = 7'h4e == _GEN_793 ? io_FromL1 : L0Memory_78; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_208 = 7'h4f == _GEN_793 ? io_FromL1 : L0Memory_79; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_209 = 7'h50 == _GEN_793 ? io_FromL1 : L0Memory_80; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_210 = 7'h51 == _GEN_793 ? io_FromL1 : L0Memory_81; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_211 = 7'h52 == _GEN_793 ? io_FromL1 : L0Memory_82; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_212 = 7'h53 == _GEN_793 ? io_FromL1 : L0Memory_83; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_213 = 7'h54 == _GEN_793 ? io_FromL1 : L0Memory_84; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_214 = 7'h55 == _GEN_793 ? io_FromL1 : L0Memory_85; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_215 = 7'h56 == _GEN_793 ? io_FromL1 : L0Memory_86; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_216 = 7'h57 == _GEN_793 ? io_FromL1 : L0Memory_87; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_217 = 7'h58 == _GEN_793 ? io_FromL1 : L0Memory_88; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_218 = 7'h59 == _GEN_793 ? io_FromL1 : L0Memory_89; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_219 = 7'h5a == _GEN_793 ? io_FromL1 : L0Memory_90; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_220 = 7'h5b == _GEN_793 ? io_FromL1 : L0Memory_91; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_221 = 7'h5c == _GEN_793 ? io_FromL1 : L0Memory_92; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_222 = 7'h5d == _GEN_793 ? io_FromL1 : L0Memory_93; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_223 = 7'h5e == _GEN_793 ? io_FromL1 : L0Memory_94; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_224 = 7'h5f == _GEN_793 ? io_FromL1 : L0Memory_95; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_225 = 7'h60 == _GEN_793 ? io_FromL1 : L0Memory_96; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_226 = 7'h61 == _GEN_793 ? io_FromL1 : L0Memory_97; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_227 = 7'h62 == _GEN_793 ? io_FromL1 : L0Memory_98; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_228 = 7'h63 == _GEN_793 ? io_FromL1 : L0Memory_99; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [5:0] _L0Index_T_2 = L0Index + 6'h1; // @[PEArray.scala 200:28]
  wire [15:0] _GEN_229 = count >= 10'h1 & count <= _T_27 ? _GEN_129 : L0Memory_0; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_230 = count >= 10'h1 & count <= _T_27 ? _GEN_130 : L0Memory_1; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_231 = count >= 10'h1 & count <= _T_27 ? _GEN_131 : L0Memory_2; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_232 = count >= 10'h1 & count <= _T_27 ? _GEN_132 : L0Memory_3; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_233 = count >= 10'h1 & count <= _T_27 ? _GEN_133 : L0Memory_4; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_234 = count >= 10'h1 & count <= _T_27 ? _GEN_134 : L0Memory_5; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_235 = count >= 10'h1 & count <= _T_27 ? _GEN_135 : L0Memory_6; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_236 = count >= 10'h1 & count <= _T_27 ? _GEN_136 : L0Memory_7; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_237 = count >= 10'h1 & count <= _T_27 ? _GEN_137 : L0Memory_8; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_238 = count >= 10'h1 & count <= _T_27 ? _GEN_138 : L0Memory_9; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_239 = count >= 10'h1 & count <= _T_27 ? _GEN_139 : L0Memory_10; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_240 = count >= 10'h1 & count <= _T_27 ? _GEN_140 : L0Memory_11; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_241 = count >= 10'h1 & count <= _T_27 ? _GEN_141 : L0Memory_12; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_242 = count >= 10'h1 & count <= _T_27 ? _GEN_142 : L0Memory_13; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_243 = count >= 10'h1 & count <= _T_27 ? _GEN_143 : L0Memory_14; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_244 = count >= 10'h1 & count <= _T_27 ? _GEN_144 : L0Memory_15; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_245 = count >= 10'h1 & count <= _T_27 ? _GEN_145 : L0Memory_16; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_246 = count >= 10'h1 & count <= _T_27 ? _GEN_146 : L0Memory_17; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_247 = count >= 10'h1 & count <= _T_27 ? _GEN_147 : L0Memory_18; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_248 = count >= 10'h1 & count <= _T_27 ? _GEN_148 : L0Memory_19; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_249 = count >= 10'h1 & count <= _T_27 ? _GEN_149 : L0Memory_20; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_250 = count >= 10'h1 & count <= _T_27 ? _GEN_150 : L0Memory_21; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_251 = count >= 10'h1 & count <= _T_27 ? _GEN_151 : L0Memory_22; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_252 = count >= 10'h1 & count <= _T_27 ? _GEN_152 : L0Memory_23; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_253 = count >= 10'h1 & count <= _T_27 ? _GEN_153 : L0Memory_24; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_254 = count >= 10'h1 & count <= _T_27 ? _GEN_154 : L0Memory_25; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_255 = count >= 10'h1 & count <= _T_27 ? _GEN_155 : L0Memory_26; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_256 = count >= 10'h1 & count <= _T_27 ? _GEN_156 : L0Memory_27; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_257 = count >= 10'h1 & count <= _T_27 ? _GEN_157 : L0Memory_28; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_258 = count >= 10'h1 & count <= _T_27 ? _GEN_158 : L0Memory_29; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_259 = count >= 10'h1 & count <= _T_27 ? _GEN_159 : L0Memory_30; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_260 = count >= 10'h1 & count <= _T_27 ? _GEN_160 : L0Memory_31; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_261 = count >= 10'h1 & count <= _T_27 ? _GEN_161 : L0Memory_32; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_262 = count >= 10'h1 & count <= _T_27 ? _GEN_162 : L0Memory_33; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_263 = count >= 10'h1 & count <= _T_27 ? _GEN_163 : L0Memory_34; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_264 = count >= 10'h1 & count <= _T_27 ? _GEN_164 : L0Memory_35; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_265 = count >= 10'h1 & count <= _T_27 ? _GEN_165 : L0Memory_36; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_266 = count >= 10'h1 & count <= _T_27 ? _GEN_166 : L0Memory_37; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_267 = count >= 10'h1 & count <= _T_27 ? _GEN_167 : L0Memory_38; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_268 = count >= 10'h1 & count <= _T_27 ? _GEN_168 : L0Memory_39; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_269 = count >= 10'h1 & count <= _T_27 ? _GEN_169 : L0Memory_40; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_270 = count >= 10'h1 & count <= _T_27 ? _GEN_170 : L0Memory_41; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_271 = count >= 10'h1 & count <= _T_27 ? _GEN_171 : L0Memory_42; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_272 = count >= 10'h1 & count <= _T_27 ? _GEN_172 : L0Memory_43; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_273 = count >= 10'h1 & count <= _T_27 ? _GEN_173 : L0Memory_44; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_274 = count >= 10'h1 & count <= _T_27 ? _GEN_174 : L0Memory_45; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_275 = count >= 10'h1 & count <= _T_27 ? _GEN_175 : L0Memory_46; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_276 = count >= 10'h1 & count <= _T_27 ? _GEN_176 : L0Memory_47; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_277 = count >= 10'h1 & count <= _T_27 ? _GEN_177 : L0Memory_48; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_278 = count >= 10'h1 & count <= _T_27 ? _GEN_178 : L0Memory_49; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_279 = count >= 10'h1 & count <= _T_27 ? _GEN_179 : L0Memory_50; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_280 = count >= 10'h1 & count <= _T_27 ? _GEN_180 : L0Memory_51; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_281 = count >= 10'h1 & count <= _T_27 ? _GEN_181 : L0Memory_52; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_282 = count >= 10'h1 & count <= _T_27 ? _GEN_182 : L0Memory_53; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_283 = count >= 10'h1 & count <= _T_27 ? _GEN_183 : L0Memory_54; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_284 = count >= 10'h1 & count <= _T_27 ? _GEN_184 : L0Memory_55; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_285 = count >= 10'h1 & count <= _T_27 ? _GEN_185 : L0Memory_56; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_286 = count >= 10'h1 & count <= _T_27 ? _GEN_186 : L0Memory_57; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_287 = count >= 10'h1 & count <= _T_27 ? _GEN_187 : L0Memory_58; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_288 = count >= 10'h1 & count <= _T_27 ? _GEN_188 : L0Memory_59; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_289 = count >= 10'h1 & count <= _T_27 ? _GEN_189 : L0Memory_60; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_290 = count >= 10'h1 & count <= _T_27 ? _GEN_190 : L0Memory_61; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_291 = count >= 10'h1 & count <= _T_27 ? _GEN_191 : L0Memory_62; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_292 = count >= 10'h1 & count <= _T_27 ? _GEN_192 : L0Memory_63; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_293 = count >= 10'h1 & count <= _T_27 ? _GEN_193 : L0Memory_64; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_294 = count >= 10'h1 & count <= _T_27 ? _GEN_194 : L0Memory_65; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_295 = count >= 10'h1 & count <= _T_27 ? _GEN_195 : L0Memory_66; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_296 = count >= 10'h1 & count <= _T_27 ? _GEN_196 : L0Memory_67; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_297 = count >= 10'h1 & count <= _T_27 ? _GEN_197 : L0Memory_68; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_298 = count >= 10'h1 & count <= _T_27 ? _GEN_198 : L0Memory_69; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_299 = count >= 10'h1 & count <= _T_27 ? _GEN_199 : L0Memory_70; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_300 = count >= 10'h1 & count <= _T_27 ? _GEN_200 : L0Memory_71; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_301 = count >= 10'h1 & count <= _T_27 ? _GEN_201 : L0Memory_72; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_302 = count >= 10'h1 & count <= _T_27 ? _GEN_202 : L0Memory_73; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_303 = count >= 10'h1 & count <= _T_27 ? _GEN_203 : L0Memory_74; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_304 = count >= 10'h1 & count <= _T_27 ? _GEN_204 : L0Memory_75; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_305 = count >= 10'h1 & count <= _T_27 ? _GEN_205 : L0Memory_76; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_306 = count >= 10'h1 & count <= _T_27 ? _GEN_206 : L0Memory_77; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_307 = count >= 10'h1 & count <= _T_27 ? _GEN_207 : L0Memory_78; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_308 = count >= 10'h1 & count <= _T_27 ? _GEN_208 : L0Memory_79; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_309 = count >= 10'h1 & count <= _T_27 ? _GEN_209 : L0Memory_80; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_310 = count >= 10'h1 & count <= _T_27 ? _GEN_210 : L0Memory_81; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_311 = count >= 10'h1 & count <= _T_27 ? _GEN_211 : L0Memory_82; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_312 = count >= 10'h1 & count <= _T_27 ? _GEN_212 : L0Memory_83; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_313 = count >= 10'h1 & count <= _T_27 ? _GEN_213 : L0Memory_84; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_314 = count >= 10'h1 & count <= _T_27 ? _GEN_214 : L0Memory_85; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_315 = count >= 10'h1 & count <= _T_27 ? _GEN_215 : L0Memory_86; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_316 = count >= 10'h1 & count <= _T_27 ? _GEN_216 : L0Memory_87; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_317 = count >= 10'h1 & count <= _T_27 ? _GEN_217 : L0Memory_88; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_318 = count >= 10'h1 & count <= _T_27 ? _GEN_218 : L0Memory_89; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_319 = count >= 10'h1 & count <= _T_27 ? _GEN_219 : L0Memory_90; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_320 = count >= 10'h1 & count <= _T_27 ? _GEN_220 : L0Memory_91; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_321 = count >= 10'h1 & count <= _T_27 ? _GEN_221 : L0Memory_92; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_322 = count >= 10'h1 & count <= _T_27 ? _GEN_222 : L0Memory_93; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_323 = count >= 10'h1 & count <= _T_27 ? _GEN_223 : L0Memory_94; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_324 = count >= 10'h1 & count <= _T_27 ? _GEN_224 : L0Memory_95; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_325 = count >= 10'h1 & count <= _T_27 ? _GEN_225 : L0Memory_96; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_326 = count >= 10'h1 & count <= _T_27 ? _GEN_226 : L0Memory_97; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_327 = count >= 10'h1 & count <= _T_27 ? _GEN_227 : L0Memory_98; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_328 = count >= 10'h1 & count <= _T_27 ? _GEN_228 : L0Memory_99; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [5:0] _GEN_329 = count >= 10'h1 & count <= _T_27 ? _L0Index_T_2 : _GEN_128; // @[PEArray.scala 198:59 PEArray.scala 200:17]
  wire [9:0] _GEN_330 = _T_24 ? 10'h0 : _GEN_127; // @[PEArray.scala 202:32 PEArray.scala 203:15]
  wire [2:0] _GEN_331 = _T_24 ? 3'h0 : state; // @[PEArray.scala 202:32 PEArray.scala 204:15 PEArray.scala 100:22]
  wire [9:0] _GEN_865 = {{4'd0}, GRU_out_width}; // @[PEArray.scala 220:19]
  wire [9:0] _GEN_0 = count % _GEN_865; // @[PEArray.scala 220:19]
  wire [5:0] _T_36 = _GEN_0[5:0]; // @[PEArray.scala 220:19]
  wire [5:0] _T_38 = GRU_out_width - 6'h1; // @[PEArray.scala 220:55]
  wire [5:0] _GEN_334 = _T_36 == _T_38 ? _L0Index_T_2 : 6'h0; // @[PEArray.scala 220:62 PEArray.scala 221:17 PEArray.scala 214:15]
  wire [5:0] _GEN_346 = _T_41 ? _GEN_334 : L0Index; // @[Conditional.scala 39:67 PEArray.scala 39:24]
  wire [9:0] _GEN_347 = _T_41 ? _GEN_330 : count; // @[Conditional.scala 39:67 PEArray.scala 101:22]
  wire [2:0] _GEN_348 = _T_41 ? _GEN_331 : state; // @[Conditional.scala 39:67 PEArray.scala 100:22]
  wire [5:0] _GEN_353 = _T_31 ? _GEN_334 : _GEN_346; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_354 = _T_31 ? _GEN_330 : _GEN_347; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_355 = _T_31 ? _GEN_331 : _GEN_348; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_356 = _T_22 ? _GEN_330 : _GEN_354; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_357 = _T_22 ? _GEN_329 : _GEN_353; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_458 = _T_22 ? _GEN_331 : _GEN_355; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_690 = _T_3 ? _GEN_118 : {{2'd0}, GRU_out_width}; // @[Conditional.scala 40:58 PEArray.scala 104:26]
  FP16MulAdder FP16MAC ( // @[PEArray.scala 72:23]
    .io_a(FP16MAC_io_a),
    .io_b(FP16MAC_io_b),
    .io_c(FP16MAC_io_c),
    .io_out(FP16MAC_io_out)
  );
  assign io_ToRightPE = mux3out_reg; // @[PEArray.scala 95:16]
  assign io_ToBelowPE = mux2out_reg; // @[PEArray.scala 94:16]
  assign FP16MAC_io_a = sel1 ? io_FromL1 : io_FromLeftPE; // @[PEArray.scala 50:14 PEArray.scala 50:23 PEArray.scala 51:24]
  assign FP16MAC_io_b = sel5 ? mux4out : _GEN_105; // @[PEArray.scala 77:13 PEArray.scala 78:18 PEArray.scala 81:18]
  assign FP16MAC_io_c = sel5 ? _GEN_105 : mux4out; // @[PEArray.scala 77:13 PEArray.scala 79:18 PEArray.scala 82:18]
  always @(posedge clock) begin
    if (reset) begin // @[PEArray.scala 39:24]
      L0Index <= 6'h0; // @[PEArray.scala 39:24]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h0; // @[PEArray.scala 159:15]
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h7; // @[PEArray.scala 181:15]
      end else begin
        L0Index <= _GEN_357;
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_0 <= _GEN_229;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_1 <= _GEN_230;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_2 <= _GEN_231;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_3 <= _GEN_232;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_4 <= _GEN_233;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_5 <= _GEN_234;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_6 <= _GEN_235;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_7 <= _GEN_236;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_8 <= _GEN_237;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_9 <= _GEN_238;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_10 <= _GEN_239;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_11 <= _GEN_240;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_12 <= _GEN_241;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_13 <= _GEN_242;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_14 <= _GEN_243;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_15 <= _GEN_244;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_16 <= _GEN_245;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_17 <= _GEN_246;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_18 <= _GEN_247;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_19 <= _GEN_248;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_20 <= _GEN_249;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_21 <= _GEN_250;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_22 <= _GEN_251;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_23 <= _GEN_252;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_24 <= _GEN_253;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_25 <= _GEN_254;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_26 <= _GEN_255;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_27 <= _GEN_256;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_28 <= _GEN_257;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_29 <= _GEN_258;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_30 <= _GEN_259;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_31 <= _GEN_260;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_32 <= _GEN_261;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_33 <= _GEN_262;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_34 <= _GEN_263;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_35 <= _GEN_264;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_36 <= _GEN_265;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_37 <= _GEN_266;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_38 <= _GEN_267;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_39 <= _GEN_268;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_40 <= _GEN_269;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_41 <= _GEN_270;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_42 <= _GEN_271;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_43 <= _GEN_272;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_44 <= _GEN_273;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_45 <= _GEN_274;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_46 <= _GEN_275;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_47 <= _GEN_276;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_48 <= _GEN_277;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_49 <= _GEN_278;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_50 <= _GEN_279;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_51 <= _GEN_280;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_52 <= _GEN_281;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_53 <= _GEN_282;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_54 <= _GEN_283;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_55 <= _GEN_284;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_56 <= _GEN_285;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_57 <= _GEN_286;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_58 <= _GEN_287;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_59 <= _GEN_288;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_60 <= _GEN_289;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_61 <= _GEN_290;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_62 <= _GEN_291;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_63 <= _GEN_292;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_64 <= _GEN_293;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_65 <= _GEN_294;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_66 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_67 <= _GEN_296;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_68 <= _GEN_297;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_69 <= _GEN_298;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_70 <= _GEN_299;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_71 <= _GEN_300;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_72 <= _GEN_301;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_73 <= _GEN_302;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_74 <= _GEN_303;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_75 <= _GEN_304;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_76 <= _GEN_305;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_77 <= _GEN_306;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_78 <= _GEN_307;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_79 <= _GEN_308;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_80 <= _GEN_309;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_81 <= _GEN_310;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_82 <= _GEN_311;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_83 <= _GEN_312;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_84 <= _GEN_313;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_85 <= _GEN_314;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_86 <= _GEN_315;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_87 <= _GEN_316;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_88 <= _GEN_317;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_89 <= _GEN_318;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_90 <= _GEN_319;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_91 <= _GEN_320;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_92 <= _GEN_321;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_93 <= _GEN_322;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_94 <= _GEN_323;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_95 <= _GEN_324;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_96 <= _GEN_325;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_97 <= _GEN_326;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_98 <= _GEN_327;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_99 <= _GEN_328;
          end
        end
      end
    end
    if (reset) begin // @[PEArray.scala 100:22]
      state <= 3'h0; // @[PEArray.scala 100:22]
    end else if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[7]) begin // @[PEArray.scala 116:57]
        state <= 3'h1;
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      if (count == 10'h33) begin // @[PEArray.scala 164:27]
        state <= 3'h0; // @[PEArray.scala 166:15]
      end
    end else if (_T_16) begin // @[Conditional.scala 39:67]
      state <= _GEN_126;
    end else begin
      state <= _GEN_458;
    end
    if (reset) begin // @[PEArray.scala 90:28]
      mux2out_reg <= 16'h0; // @[PEArray.scala 90:28]
    end else begin
      mux2out_reg <= MAC_out; // @[PEArray.scala 90:28]
    end
    if (reset) begin // @[PEArray.scala 91:28]
      mux3out_reg <= 16'h0; // @[PEArray.scala 91:28]
    end else if (sel3) begin // @[PEArray.scala 56:14]
      mux3out_reg <= MAC_out; // @[PEArray.scala 56:23]
    end else if (sel1) begin // @[PEArray.scala 50:14]
      mux3out_reg <= io_FromL1; // @[PEArray.scala 50:23]
    end else begin
      mux3out_reg <= io_FromLeftPE; // @[PEArray.scala 51:24]
    end
    if (reset) begin // @[PEArray.scala 101:22]
      count <= 10'h0; // @[PEArray.scala 101:22]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        if (count == 10'h33) begin // @[PEArray.scala 164:27]
          count <= 10'h0; // @[PEArray.scala 165:15]
        end else begin
          count <= _GEN_120;
        end
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        count <= _GEN_125;
      end else begin
        count <= _GEN_356;
      end
    end
    GRU_out_width <= _GEN_690[5:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  L0Index = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  L0Memory_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  L0Memory_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  L0Memory_2 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  L0Memory_3 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  L0Memory_4 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  L0Memory_5 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  L0Memory_6 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  L0Memory_7 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  L0Memory_8 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  L0Memory_9 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  L0Memory_10 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  L0Memory_11 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  L0Memory_12 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  L0Memory_13 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  L0Memory_14 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  L0Memory_15 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  L0Memory_16 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  L0Memory_17 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  L0Memory_18 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  L0Memory_19 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  L0Memory_20 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  L0Memory_21 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  L0Memory_22 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  L0Memory_23 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  L0Memory_24 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  L0Memory_25 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  L0Memory_26 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  L0Memory_27 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  L0Memory_28 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  L0Memory_29 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  L0Memory_30 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  L0Memory_31 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  L0Memory_32 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  L0Memory_33 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  L0Memory_34 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  L0Memory_35 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  L0Memory_36 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  L0Memory_37 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  L0Memory_38 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  L0Memory_39 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  L0Memory_40 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  L0Memory_41 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  L0Memory_42 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  L0Memory_43 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  L0Memory_44 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  L0Memory_45 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  L0Memory_46 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  L0Memory_47 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  L0Memory_48 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  L0Memory_49 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  L0Memory_50 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  L0Memory_51 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  L0Memory_52 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  L0Memory_53 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  L0Memory_54 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  L0Memory_55 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  L0Memory_56 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  L0Memory_57 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  L0Memory_58 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  L0Memory_59 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  L0Memory_60 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  L0Memory_61 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  L0Memory_62 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  L0Memory_63 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  L0Memory_64 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  L0Memory_65 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  L0Memory_66 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  L0Memory_67 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  L0Memory_68 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  L0Memory_69 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  L0Memory_70 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  L0Memory_71 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  L0Memory_72 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  L0Memory_73 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  L0Memory_74 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  L0Memory_75 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  L0Memory_76 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  L0Memory_77 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  L0Memory_78 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  L0Memory_79 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  L0Memory_80 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  L0Memory_81 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  L0Memory_82 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  L0Memory_83 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  L0Memory_84 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  L0Memory_85 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  L0Memory_86 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  L0Memory_87 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  L0Memory_88 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  L0Memory_89 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  L0Memory_90 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  L0Memory_91 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  L0Memory_92 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  L0Memory_93 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  L0Memory_94 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  L0Memory_95 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  L0Memory_96 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  L0Memory_97 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  L0Memory_98 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  L0Memory_99 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  state = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  mux2out_reg = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  mux3out_reg = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  count = _RAND_104[9:0];
  _RAND_105 = {1{`RANDOM}};
  GRU_out_width = _RAND_105[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PE_13(
  input         clock,
  input         reset,
  input  [15:0] io_FromAbovePE,
  input  [15:0] io_FromLeftPE,
  input  [15:0] io_FromL1,
  input  [11:0] io_control_signal_mask,
  output [15:0] io_ToRightPE,
  output [15:0] io_ToBelowPE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] FP16MAC_io_a; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_b; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_c; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_out; // @[PEArray.scala 72:23]
  reg [5:0] L0Index; // @[PEArray.scala 39:24]
  reg [15:0] L0Memory_0; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_1; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_2; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_3; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_4; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_5; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_6; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_7; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_8; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_9; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_10; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_11; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_12; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_13; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_14; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_15; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_16; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_17; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_18; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_19; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_20; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_21; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_22; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_23; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_24; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_25; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_26; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_27; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_28; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_29; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_30; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_31; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_32; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_33; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_34; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_35; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_36; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_37; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_38; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_39; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_40; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_41; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_42; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_43; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_44; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_45; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_46; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_47; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_48; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_49; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_50; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_51; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_52; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_53; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_54; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_55; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_56; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_57; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_58; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_59; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_60; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_61; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_62; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_63; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_64; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_65; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_66; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_67; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_68; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_69; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_70; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_71; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_72; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_73; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_74; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_75; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_76; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_77; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_78; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_79; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_80; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_81; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_82; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_83; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_84; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_85; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_86; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_87; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_88; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_89; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_90; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_91; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_92; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_93; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_94; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_95; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_96; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_97; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_98; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_99; // @[PEArray.scala 40:21]
  reg [2:0] state; // @[PEArray.scala 100:22]
  wire  _T_3 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_12 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_16 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_22 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_31 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_41 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_342 = _T_41 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 231:12 PEArray.scala 32:8]
  wire  _GEN_349 = _T_31 ? 1'h0 : _GEN_342; // @[Conditional.scala 39:67 PEArray.scala 208:12]
  wire  _GEN_459 = _T_22 | _GEN_349; // @[Conditional.scala 39:67 PEArray.scala 32:8]
  wire  _GEN_463 = _T_16 ? 1'h0 : _GEN_459; // @[Conditional.scala 39:67]
  wire  _GEN_572 = _T_12 | _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 149:12]
  wire  sel1 = _T_3 | _GEN_572; // @[Conditional.scala 40:58 PEArray.scala 108:12]
  wire [15:0] MAC_out = FP16MAC_io_out; // @[PEArray.scala 47:21 PEArray.scala 85:11]
  wire  _GEN_465 = _T_16 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 177:12]
  wire  _GEN_580 = _T_12 | _GEN_465; // @[Conditional.scala 39:67 PEArray.scala 34:8]
  wire  sel3 = _T_3 | _GEN_580; // @[Conditional.scala 40:58 PEArray.scala 110:12]
  wire [1:0] _GEN_344 = _T_41 ? 2'h2 : 2'h0; // @[Conditional.scala 39:67 PEArray.scala 233:12 PEArray.scala 35:8]
  wire [1:0] _GEN_351 = _T_31 ? 2'h2 : _GEN_344; // @[Conditional.scala 39:67 PEArray.scala 210:12]
  wire [1:0] _GEN_461 = _T_22 ? 2'h0 : _GEN_351; // @[Conditional.scala 39:67 PEArray.scala 35:8]
  wire [1:0] _GEN_466 = _T_16 ? 2'h0 : _GEN_461; // @[Conditional.scala 39:67 PEArray.scala 178:12]
  wire [1:0] _GEN_574 = _T_12 ? 2'h1 : _GEN_466; // @[Conditional.scala 39:67]
  wire [1:0] sel4 = _T_3 ? 2'h0 : _GEN_574; // @[Conditional.scala 40:58 PEArray.scala 111:12]
  wire [15:0] _GEN_3 = sel4 == 2'h2 ? io_FromL1 : 16'h0; // @[PEArray.scala 65:28 PEArray.scala 66:15 PEArray.scala 69:15]
  wire [15:0] _GEN_4 = sel4 == 2'h1 ? io_FromAbovePE : _GEN_3; // @[PEArray.scala 62:28 PEArray.scala 63:15]
  wire [15:0] mux4out = sel4 == 2'h0 ? 16'h0 : _GEN_4; // @[PEArray.scala 59:22 PEArray.scala 60:13]
  wire [15:0] _GEN_7 = 6'h1 == L0Index ? L0Memory_1 : L0Memory_0; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_8 = 6'h2 == L0Index ? L0Memory_2 : _GEN_7; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_9 = 6'h3 == L0Index ? L0Memory_3 : _GEN_8; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_10 = 6'h4 == L0Index ? L0Memory_4 : _GEN_9; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_11 = 6'h5 == L0Index ? L0Memory_5 : _GEN_10; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_12 = 6'h6 == L0Index ? L0Memory_6 : _GEN_11; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_13 = 6'h7 == L0Index ? L0Memory_7 : _GEN_12; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_14 = 6'h8 == L0Index ? L0Memory_8 : _GEN_13; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_15 = 6'h9 == L0Index ? L0Memory_9 : _GEN_14; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_16 = 6'ha == L0Index ? L0Memory_10 : _GEN_15; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_17 = 6'hb == L0Index ? L0Memory_11 : _GEN_16; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_18 = 6'hc == L0Index ? L0Memory_12 : _GEN_17; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_19 = 6'hd == L0Index ? L0Memory_13 : _GEN_18; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_20 = 6'he == L0Index ? L0Memory_14 : _GEN_19; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_21 = 6'hf == L0Index ? L0Memory_15 : _GEN_20; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_22 = 6'h10 == L0Index ? L0Memory_16 : _GEN_21; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_23 = 6'h11 == L0Index ? L0Memory_17 : _GEN_22; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_24 = 6'h12 == L0Index ? L0Memory_18 : _GEN_23; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_25 = 6'h13 == L0Index ? L0Memory_19 : _GEN_24; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_26 = 6'h14 == L0Index ? L0Memory_20 : _GEN_25; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_27 = 6'h15 == L0Index ? L0Memory_21 : _GEN_26; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_28 = 6'h16 == L0Index ? L0Memory_22 : _GEN_27; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_29 = 6'h17 == L0Index ? L0Memory_23 : _GEN_28; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_30 = 6'h18 == L0Index ? L0Memory_24 : _GEN_29; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_31 = 6'h19 == L0Index ? L0Memory_25 : _GEN_30; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_32 = 6'h1a == L0Index ? L0Memory_26 : _GEN_31; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_33 = 6'h1b == L0Index ? L0Memory_27 : _GEN_32; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_34 = 6'h1c == L0Index ? L0Memory_28 : _GEN_33; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_35 = 6'h1d == L0Index ? L0Memory_29 : _GEN_34; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_36 = 6'h1e == L0Index ? L0Memory_30 : _GEN_35; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_37 = 6'h1f == L0Index ? L0Memory_31 : _GEN_36; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_38 = 6'h20 == L0Index ? L0Memory_32 : _GEN_37; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_39 = 6'h21 == L0Index ? L0Memory_33 : _GEN_38; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_40 = 6'h22 == L0Index ? L0Memory_34 : _GEN_39; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_41 = 6'h23 == L0Index ? L0Memory_35 : _GEN_40; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_42 = 6'h24 == L0Index ? L0Memory_36 : _GEN_41; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_43 = 6'h25 == L0Index ? L0Memory_37 : _GEN_42; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_44 = 6'h26 == L0Index ? L0Memory_38 : _GEN_43; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_45 = 6'h27 == L0Index ? L0Memory_39 : _GEN_44; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_46 = 6'h28 == L0Index ? L0Memory_40 : _GEN_45; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_47 = 6'h29 == L0Index ? L0Memory_41 : _GEN_46; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_48 = 6'h2a == L0Index ? L0Memory_42 : _GEN_47; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_49 = 6'h2b == L0Index ? L0Memory_43 : _GEN_48; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_50 = 6'h2c == L0Index ? L0Memory_44 : _GEN_49; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_51 = 6'h2d == L0Index ? L0Memory_45 : _GEN_50; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_52 = 6'h2e == L0Index ? L0Memory_46 : _GEN_51; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_53 = 6'h2f == L0Index ? L0Memory_47 : _GEN_52; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_54 = 6'h30 == L0Index ? L0Memory_48 : _GEN_53; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_55 = 6'h31 == L0Index ? L0Memory_49 : _GEN_54; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_56 = 6'h32 == L0Index ? L0Memory_50 : _GEN_55; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_57 = 6'h33 == L0Index ? L0Memory_51 : _GEN_56; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_58 = 6'h34 == L0Index ? L0Memory_52 : _GEN_57; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_59 = 6'h35 == L0Index ? L0Memory_53 : _GEN_58; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_60 = 6'h36 == L0Index ? L0Memory_54 : _GEN_59; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_61 = 6'h37 == L0Index ? L0Memory_55 : _GEN_60; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_62 = 6'h38 == L0Index ? L0Memory_56 : _GEN_61; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_63 = 6'h39 == L0Index ? L0Memory_57 : _GEN_62; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_64 = 6'h3a == L0Index ? L0Memory_58 : _GEN_63; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_65 = 6'h3b == L0Index ? L0Memory_59 : _GEN_64; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_66 = 6'h3c == L0Index ? L0Memory_60 : _GEN_65; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_67 = 6'h3d == L0Index ? L0Memory_61 : _GEN_66; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_68 = 6'h3e == L0Index ? L0Memory_62 : _GEN_67; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_69 = 6'h3f == L0Index ? L0Memory_63 : _GEN_68; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [6:0] _GEN_793 = {{1'd0}, L0Index}; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_70 = 7'h40 == _GEN_793 ? L0Memory_64 : _GEN_69; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_71 = 7'h41 == _GEN_793 ? L0Memory_65 : _GEN_70; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_72 = 7'h42 == _GEN_793 ? L0Memory_66 : _GEN_71; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_73 = 7'h43 == _GEN_793 ? L0Memory_67 : _GEN_72; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_74 = 7'h44 == _GEN_793 ? L0Memory_68 : _GEN_73; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_75 = 7'h45 == _GEN_793 ? L0Memory_69 : _GEN_74; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_76 = 7'h46 == _GEN_793 ? L0Memory_70 : _GEN_75; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_77 = 7'h47 == _GEN_793 ? L0Memory_71 : _GEN_76; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_78 = 7'h48 == _GEN_793 ? L0Memory_72 : _GEN_77; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_79 = 7'h49 == _GEN_793 ? L0Memory_73 : _GEN_78; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_80 = 7'h4a == _GEN_793 ? L0Memory_74 : _GEN_79; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_81 = 7'h4b == _GEN_793 ? L0Memory_75 : _GEN_80; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_82 = 7'h4c == _GEN_793 ? L0Memory_76 : _GEN_81; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_83 = 7'h4d == _GEN_793 ? L0Memory_77 : _GEN_82; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_84 = 7'h4e == _GEN_793 ? L0Memory_78 : _GEN_83; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_85 = 7'h4f == _GEN_793 ? L0Memory_79 : _GEN_84; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_86 = 7'h50 == _GEN_793 ? L0Memory_80 : _GEN_85; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_87 = 7'h51 == _GEN_793 ? L0Memory_81 : _GEN_86; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_88 = 7'h52 == _GEN_793 ? L0Memory_82 : _GEN_87; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_89 = 7'h53 == _GEN_793 ? L0Memory_83 : _GEN_88; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_90 = 7'h54 == _GEN_793 ? L0Memory_84 : _GEN_89; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_91 = 7'h55 == _GEN_793 ? L0Memory_85 : _GEN_90; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_92 = 7'h56 == _GEN_793 ? L0Memory_86 : _GEN_91; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_93 = 7'h57 == _GEN_793 ? L0Memory_87 : _GEN_92; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_94 = 7'h58 == _GEN_793 ? L0Memory_88 : _GEN_93; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_95 = 7'h59 == _GEN_793 ? L0Memory_89 : _GEN_94; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_96 = 7'h5a == _GEN_793 ? L0Memory_90 : _GEN_95; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_97 = 7'h5b == _GEN_793 ? L0Memory_91 : _GEN_96; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_98 = 7'h5c == _GEN_793 ? L0Memory_92 : _GEN_97; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_99 = 7'h5d == _GEN_793 ? L0Memory_93 : _GEN_98; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_100 = 7'h5e == _GEN_793 ? L0Memory_94 : _GEN_99; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_101 = 7'h5f == _GEN_793 ? L0Memory_95 : _GEN_100; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_102 = 7'h60 == _GEN_793 ? L0Memory_96 : _GEN_101; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_103 = 7'h61 == _GEN_793 ? L0Memory_97 : _GEN_102; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_104 = 7'h62 == _GEN_793 ? L0Memory_98 : _GEN_103; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_105 = 7'h63 == _GEN_793 ? L0Memory_99 : _GEN_104; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire  _GEN_575 = _T_12 ? 1'h0 : _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 157:12]
  wire  sel5 = _T_3 ? 1'h0 : _GEN_575; // @[Conditional.scala 40:58 PEArray.scala 112:12]
  reg [15:0] mux2out_reg; // @[PEArray.scala 90:28]
  reg [15:0] mux3out_reg; // @[PEArray.scala 91:28]
  reg [9:0] count; // @[PEArray.scala 101:22]
  reg [5:0] GRU_out_width; // @[PEArray.scala 104:26]
  wire [7:0] _GEN_118 = io_control_signal_mask[7] ? 8'h0 : {{2'd0}, GRU_out_width}; // @[PEArray.scala 116:57 PEArray.scala 145:23 PEArray.scala 104:26]
  wire [9:0] _count_T_1 = count + 10'h1; // @[PEArray.scala 162:24]
  wire [9:0] _GEN_120 = count != 10'h33 ? _count_T_1 : count; // @[PEArray.scala 161:27 PEArray.scala 162:15 PEArray.scala 101:22]
  wire [9:0] _GEN_124 = count != 10'h188 ? _count_T_1 : count; // @[PEArray.scala 183:28 PEArray.scala 184:15 PEArray.scala 101:22]
  wire [9:0] _GEN_125 = count == 10'h188 ? 10'h0 : _GEN_124; // @[PEArray.scala 186:28 PEArray.scala 187:15]
  wire [2:0] _GEN_126 = count == 10'h188 ? 3'h0 : state; // @[PEArray.scala 186:28 PEArray.scala 188:15 PEArray.scala 100:22]
  wire [9:0] _GEN_127 = count != 10'h0 ? _count_T_1 : count; // @[PEArray.scala 192:32 PEArray.scala 193:15 PEArray.scala 101:22]
  wire  _T_24 = count == 10'h0; // @[PEArray.scala 195:18]
  wire [5:0] _GEN_128 = count == 10'h0 ? 6'h0 : L0Index; // @[PEArray.scala 195:26 PEArray.scala 196:17 PEArray.scala 39:24]
  wire [9:0] _T_27 = 10'h0 - 10'h1; // @[PEArray.scala 198:51]
  wire [15:0] _GEN_129 = 6'h0 == L0Index ? io_FromL1 : L0Memory_0; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_130 = 6'h1 == L0Index ? io_FromL1 : L0Memory_1; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_131 = 6'h2 == L0Index ? io_FromL1 : L0Memory_2; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_132 = 6'h3 == L0Index ? io_FromL1 : L0Memory_3; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_133 = 6'h4 == L0Index ? io_FromL1 : L0Memory_4; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_134 = 6'h5 == L0Index ? io_FromL1 : L0Memory_5; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_135 = 6'h6 == L0Index ? io_FromL1 : L0Memory_6; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_136 = 6'h7 == L0Index ? io_FromL1 : L0Memory_7; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_137 = 6'h8 == L0Index ? io_FromL1 : L0Memory_8; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_138 = 6'h9 == L0Index ? io_FromL1 : L0Memory_9; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_139 = 6'ha == L0Index ? io_FromL1 : L0Memory_10; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_140 = 6'hb == L0Index ? io_FromL1 : L0Memory_11; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_141 = 6'hc == L0Index ? io_FromL1 : L0Memory_12; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_142 = 6'hd == L0Index ? io_FromL1 : L0Memory_13; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_143 = 6'he == L0Index ? io_FromL1 : L0Memory_14; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_144 = 6'hf == L0Index ? io_FromL1 : L0Memory_15; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_145 = 6'h10 == L0Index ? io_FromL1 : L0Memory_16; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_146 = 6'h11 == L0Index ? io_FromL1 : L0Memory_17; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_147 = 6'h12 == L0Index ? io_FromL1 : L0Memory_18; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_148 = 6'h13 == L0Index ? io_FromL1 : L0Memory_19; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_149 = 6'h14 == L0Index ? io_FromL1 : L0Memory_20; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_150 = 6'h15 == L0Index ? io_FromL1 : L0Memory_21; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_151 = 6'h16 == L0Index ? io_FromL1 : L0Memory_22; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_152 = 6'h17 == L0Index ? io_FromL1 : L0Memory_23; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_153 = 6'h18 == L0Index ? io_FromL1 : L0Memory_24; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_154 = 6'h19 == L0Index ? io_FromL1 : L0Memory_25; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_155 = 6'h1a == L0Index ? io_FromL1 : L0Memory_26; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_156 = 6'h1b == L0Index ? io_FromL1 : L0Memory_27; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_157 = 6'h1c == L0Index ? io_FromL1 : L0Memory_28; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_158 = 6'h1d == L0Index ? io_FromL1 : L0Memory_29; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_159 = 6'h1e == L0Index ? io_FromL1 : L0Memory_30; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_160 = 6'h1f == L0Index ? io_FromL1 : L0Memory_31; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_161 = 6'h20 == L0Index ? io_FromL1 : L0Memory_32; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_162 = 6'h21 == L0Index ? io_FromL1 : L0Memory_33; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_163 = 6'h22 == L0Index ? io_FromL1 : L0Memory_34; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_164 = 6'h23 == L0Index ? io_FromL1 : L0Memory_35; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_165 = 6'h24 == L0Index ? io_FromL1 : L0Memory_36; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_166 = 6'h25 == L0Index ? io_FromL1 : L0Memory_37; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_167 = 6'h26 == L0Index ? io_FromL1 : L0Memory_38; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_168 = 6'h27 == L0Index ? io_FromL1 : L0Memory_39; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_169 = 6'h28 == L0Index ? io_FromL1 : L0Memory_40; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_170 = 6'h29 == L0Index ? io_FromL1 : L0Memory_41; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_171 = 6'h2a == L0Index ? io_FromL1 : L0Memory_42; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_172 = 6'h2b == L0Index ? io_FromL1 : L0Memory_43; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_173 = 6'h2c == L0Index ? io_FromL1 : L0Memory_44; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_174 = 6'h2d == L0Index ? io_FromL1 : L0Memory_45; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_175 = 6'h2e == L0Index ? io_FromL1 : L0Memory_46; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_176 = 6'h2f == L0Index ? io_FromL1 : L0Memory_47; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_177 = 6'h30 == L0Index ? io_FromL1 : L0Memory_48; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_178 = 6'h31 == L0Index ? io_FromL1 : L0Memory_49; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_179 = 6'h32 == L0Index ? io_FromL1 : L0Memory_50; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_180 = 6'h33 == L0Index ? io_FromL1 : L0Memory_51; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_181 = 6'h34 == L0Index ? io_FromL1 : L0Memory_52; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_182 = 6'h35 == L0Index ? io_FromL1 : L0Memory_53; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_183 = 6'h36 == L0Index ? io_FromL1 : L0Memory_54; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_184 = 6'h37 == L0Index ? io_FromL1 : L0Memory_55; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_185 = 6'h38 == L0Index ? io_FromL1 : L0Memory_56; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_186 = 6'h39 == L0Index ? io_FromL1 : L0Memory_57; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_187 = 6'h3a == L0Index ? io_FromL1 : L0Memory_58; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_188 = 6'h3b == L0Index ? io_FromL1 : L0Memory_59; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_189 = 6'h3c == L0Index ? io_FromL1 : L0Memory_60; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_190 = 6'h3d == L0Index ? io_FromL1 : L0Memory_61; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_191 = 6'h3e == L0Index ? io_FromL1 : L0Memory_62; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_192 = 6'h3f == L0Index ? io_FromL1 : L0Memory_63; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_193 = 7'h40 == _GEN_793 ? io_FromL1 : L0Memory_64; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_194 = 7'h41 == _GEN_793 ? io_FromL1 : L0Memory_65; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_195 = 7'h42 == _GEN_793 ? io_FromL1 : L0Memory_66; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_196 = 7'h43 == _GEN_793 ? io_FromL1 : L0Memory_67; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_197 = 7'h44 == _GEN_793 ? io_FromL1 : L0Memory_68; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_198 = 7'h45 == _GEN_793 ? io_FromL1 : L0Memory_69; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_199 = 7'h46 == _GEN_793 ? io_FromL1 : L0Memory_70; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_200 = 7'h47 == _GEN_793 ? io_FromL1 : L0Memory_71; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_201 = 7'h48 == _GEN_793 ? io_FromL1 : L0Memory_72; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_202 = 7'h49 == _GEN_793 ? io_FromL1 : L0Memory_73; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_203 = 7'h4a == _GEN_793 ? io_FromL1 : L0Memory_74; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_204 = 7'h4b == _GEN_793 ? io_FromL1 : L0Memory_75; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_205 = 7'h4c == _GEN_793 ? io_FromL1 : L0Memory_76; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_206 = 7'h4d == _GEN_793 ? io_FromL1 : L0Memory_77; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_207 = 7'h4e == _GEN_793 ? io_FromL1 : L0Memory_78; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_208 = 7'h4f == _GEN_793 ? io_FromL1 : L0Memory_79; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_209 = 7'h50 == _GEN_793 ? io_FromL1 : L0Memory_80; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_210 = 7'h51 == _GEN_793 ? io_FromL1 : L0Memory_81; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_211 = 7'h52 == _GEN_793 ? io_FromL1 : L0Memory_82; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_212 = 7'h53 == _GEN_793 ? io_FromL1 : L0Memory_83; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_213 = 7'h54 == _GEN_793 ? io_FromL1 : L0Memory_84; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_214 = 7'h55 == _GEN_793 ? io_FromL1 : L0Memory_85; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_215 = 7'h56 == _GEN_793 ? io_FromL1 : L0Memory_86; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_216 = 7'h57 == _GEN_793 ? io_FromL1 : L0Memory_87; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_217 = 7'h58 == _GEN_793 ? io_FromL1 : L0Memory_88; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_218 = 7'h59 == _GEN_793 ? io_FromL1 : L0Memory_89; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_219 = 7'h5a == _GEN_793 ? io_FromL1 : L0Memory_90; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_220 = 7'h5b == _GEN_793 ? io_FromL1 : L0Memory_91; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_221 = 7'h5c == _GEN_793 ? io_FromL1 : L0Memory_92; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_222 = 7'h5d == _GEN_793 ? io_FromL1 : L0Memory_93; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_223 = 7'h5e == _GEN_793 ? io_FromL1 : L0Memory_94; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_224 = 7'h5f == _GEN_793 ? io_FromL1 : L0Memory_95; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_225 = 7'h60 == _GEN_793 ? io_FromL1 : L0Memory_96; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_226 = 7'h61 == _GEN_793 ? io_FromL1 : L0Memory_97; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_227 = 7'h62 == _GEN_793 ? io_FromL1 : L0Memory_98; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_228 = 7'h63 == _GEN_793 ? io_FromL1 : L0Memory_99; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [5:0] _L0Index_T_2 = L0Index + 6'h1; // @[PEArray.scala 200:28]
  wire [15:0] _GEN_229 = count >= 10'h1 & count <= _T_27 ? _GEN_129 : L0Memory_0; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_230 = count >= 10'h1 & count <= _T_27 ? _GEN_130 : L0Memory_1; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_231 = count >= 10'h1 & count <= _T_27 ? _GEN_131 : L0Memory_2; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_232 = count >= 10'h1 & count <= _T_27 ? _GEN_132 : L0Memory_3; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_233 = count >= 10'h1 & count <= _T_27 ? _GEN_133 : L0Memory_4; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_234 = count >= 10'h1 & count <= _T_27 ? _GEN_134 : L0Memory_5; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_235 = count >= 10'h1 & count <= _T_27 ? _GEN_135 : L0Memory_6; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_236 = count >= 10'h1 & count <= _T_27 ? _GEN_136 : L0Memory_7; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_237 = count >= 10'h1 & count <= _T_27 ? _GEN_137 : L0Memory_8; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_238 = count >= 10'h1 & count <= _T_27 ? _GEN_138 : L0Memory_9; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_239 = count >= 10'h1 & count <= _T_27 ? _GEN_139 : L0Memory_10; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_240 = count >= 10'h1 & count <= _T_27 ? _GEN_140 : L0Memory_11; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_241 = count >= 10'h1 & count <= _T_27 ? _GEN_141 : L0Memory_12; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_242 = count >= 10'h1 & count <= _T_27 ? _GEN_142 : L0Memory_13; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_243 = count >= 10'h1 & count <= _T_27 ? _GEN_143 : L0Memory_14; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_244 = count >= 10'h1 & count <= _T_27 ? _GEN_144 : L0Memory_15; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_245 = count >= 10'h1 & count <= _T_27 ? _GEN_145 : L0Memory_16; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_246 = count >= 10'h1 & count <= _T_27 ? _GEN_146 : L0Memory_17; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_247 = count >= 10'h1 & count <= _T_27 ? _GEN_147 : L0Memory_18; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_248 = count >= 10'h1 & count <= _T_27 ? _GEN_148 : L0Memory_19; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_249 = count >= 10'h1 & count <= _T_27 ? _GEN_149 : L0Memory_20; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_250 = count >= 10'h1 & count <= _T_27 ? _GEN_150 : L0Memory_21; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_251 = count >= 10'h1 & count <= _T_27 ? _GEN_151 : L0Memory_22; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_252 = count >= 10'h1 & count <= _T_27 ? _GEN_152 : L0Memory_23; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_253 = count >= 10'h1 & count <= _T_27 ? _GEN_153 : L0Memory_24; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_254 = count >= 10'h1 & count <= _T_27 ? _GEN_154 : L0Memory_25; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_255 = count >= 10'h1 & count <= _T_27 ? _GEN_155 : L0Memory_26; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_256 = count >= 10'h1 & count <= _T_27 ? _GEN_156 : L0Memory_27; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_257 = count >= 10'h1 & count <= _T_27 ? _GEN_157 : L0Memory_28; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_258 = count >= 10'h1 & count <= _T_27 ? _GEN_158 : L0Memory_29; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_259 = count >= 10'h1 & count <= _T_27 ? _GEN_159 : L0Memory_30; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_260 = count >= 10'h1 & count <= _T_27 ? _GEN_160 : L0Memory_31; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_261 = count >= 10'h1 & count <= _T_27 ? _GEN_161 : L0Memory_32; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_262 = count >= 10'h1 & count <= _T_27 ? _GEN_162 : L0Memory_33; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_263 = count >= 10'h1 & count <= _T_27 ? _GEN_163 : L0Memory_34; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_264 = count >= 10'h1 & count <= _T_27 ? _GEN_164 : L0Memory_35; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_265 = count >= 10'h1 & count <= _T_27 ? _GEN_165 : L0Memory_36; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_266 = count >= 10'h1 & count <= _T_27 ? _GEN_166 : L0Memory_37; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_267 = count >= 10'h1 & count <= _T_27 ? _GEN_167 : L0Memory_38; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_268 = count >= 10'h1 & count <= _T_27 ? _GEN_168 : L0Memory_39; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_269 = count >= 10'h1 & count <= _T_27 ? _GEN_169 : L0Memory_40; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_270 = count >= 10'h1 & count <= _T_27 ? _GEN_170 : L0Memory_41; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_271 = count >= 10'h1 & count <= _T_27 ? _GEN_171 : L0Memory_42; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_272 = count >= 10'h1 & count <= _T_27 ? _GEN_172 : L0Memory_43; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_273 = count >= 10'h1 & count <= _T_27 ? _GEN_173 : L0Memory_44; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_274 = count >= 10'h1 & count <= _T_27 ? _GEN_174 : L0Memory_45; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_275 = count >= 10'h1 & count <= _T_27 ? _GEN_175 : L0Memory_46; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_276 = count >= 10'h1 & count <= _T_27 ? _GEN_176 : L0Memory_47; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_277 = count >= 10'h1 & count <= _T_27 ? _GEN_177 : L0Memory_48; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_278 = count >= 10'h1 & count <= _T_27 ? _GEN_178 : L0Memory_49; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_279 = count >= 10'h1 & count <= _T_27 ? _GEN_179 : L0Memory_50; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_280 = count >= 10'h1 & count <= _T_27 ? _GEN_180 : L0Memory_51; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_281 = count >= 10'h1 & count <= _T_27 ? _GEN_181 : L0Memory_52; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_282 = count >= 10'h1 & count <= _T_27 ? _GEN_182 : L0Memory_53; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_283 = count >= 10'h1 & count <= _T_27 ? _GEN_183 : L0Memory_54; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_284 = count >= 10'h1 & count <= _T_27 ? _GEN_184 : L0Memory_55; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_285 = count >= 10'h1 & count <= _T_27 ? _GEN_185 : L0Memory_56; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_286 = count >= 10'h1 & count <= _T_27 ? _GEN_186 : L0Memory_57; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_287 = count >= 10'h1 & count <= _T_27 ? _GEN_187 : L0Memory_58; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_288 = count >= 10'h1 & count <= _T_27 ? _GEN_188 : L0Memory_59; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_289 = count >= 10'h1 & count <= _T_27 ? _GEN_189 : L0Memory_60; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_290 = count >= 10'h1 & count <= _T_27 ? _GEN_190 : L0Memory_61; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_291 = count >= 10'h1 & count <= _T_27 ? _GEN_191 : L0Memory_62; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_292 = count >= 10'h1 & count <= _T_27 ? _GEN_192 : L0Memory_63; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_293 = count >= 10'h1 & count <= _T_27 ? _GEN_193 : L0Memory_64; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_294 = count >= 10'h1 & count <= _T_27 ? _GEN_194 : L0Memory_65; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_295 = count >= 10'h1 & count <= _T_27 ? _GEN_195 : L0Memory_66; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_296 = count >= 10'h1 & count <= _T_27 ? _GEN_196 : L0Memory_67; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_297 = count >= 10'h1 & count <= _T_27 ? _GEN_197 : L0Memory_68; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_298 = count >= 10'h1 & count <= _T_27 ? _GEN_198 : L0Memory_69; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_299 = count >= 10'h1 & count <= _T_27 ? _GEN_199 : L0Memory_70; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_300 = count >= 10'h1 & count <= _T_27 ? _GEN_200 : L0Memory_71; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_301 = count >= 10'h1 & count <= _T_27 ? _GEN_201 : L0Memory_72; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_302 = count >= 10'h1 & count <= _T_27 ? _GEN_202 : L0Memory_73; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_303 = count >= 10'h1 & count <= _T_27 ? _GEN_203 : L0Memory_74; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_304 = count >= 10'h1 & count <= _T_27 ? _GEN_204 : L0Memory_75; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_305 = count >= 10'h1 & count <= _T_27 ? _GEN_205 : L0Memory_76; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_306 = count >= 10'h1 & count <= _T_27 ? _GEN_206 : L0Memory_77; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_307 = count >= 10'h1 & count <= _T_27 ? _GEN_207 : L0Memory_78; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_308 = count >= 10'h1 & count <= _T_27 ? _GEN_208 : L0Memory_79; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_309 = count >= 10'h1 & count <= _T_27 ? _GEN_209 : L0Memory_80; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_310 = count >= 10'h1 & count <= _T_27 ? _GEN_210 : L0Memory_81; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_311 = count >= 10'h1 & count <= _T_27 ? _GEN_211 : L0Memory_82; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_312 = count >= 10'h1 & count <= _T_27 ? _GEN_212 : L0Memory_83; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_313 = count >= 10'h1 & count <= _T_27 ? _GEN_213 : L0Memory_84; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_314 = count >= 10'h1 & count <= _T_27 ? _GEN_214 : L0Memory_85; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_315 = count >= 10'h1 & count <= _T_27 ? _GEN_215 : L0Memory_86; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_316 = count >= 10'h1 & count <= _T_27 ? _GEN_216 : L0Memory_87; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_317 = count >= 10'h1 & count <= _T_27 ? _GEN_217 : L0Memory_88; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_318 = count >= 10'h1 & count <= _T_27 ? _GEN_218 : L0Memory_89; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_319 = count >= 10'h1 & count <= _T_27 ? _GEN_219 : L0Memory_90; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_320 = count >= 10'h1 & count <= _T_27 ? _GEN_220 : L0Memory_91; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_321 = count >= 10'h1 & count <= _T_27 ? _GEN_221 : L0Memory_92; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_322 = count >= 10'h1 & count <= _T_27 ? _GEN_222 : L0Memory_93; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_323 = count >= 10'h1 & count <= _T_27 ? _GEN_223 : L0Memory_94; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_324 = count >= 10'h1 & count <= _T_27 ? _GEN_224 : L0Memory_95; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_325 = count >= 10'h1 & count <= _T_27 ? _GEN_225 : L0Memory_96; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_326 = count >= 10'h1 & count <= _T_27 ? _GEN_226 : L0Memory_97; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_327 = count >= 10'h1 & count <= _T_27 ? _GEN_227 : L0Memory_98; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_328 = count >= 10'h1 & count <= _T_27 ? _GEN_228 : L0Memory_99; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [5:0] _GEN_329 = count >= 10'h1 & count <= _T_27 ? _L0Index_T_2 : _GEN_128; // @[PEArray.scala 198:59 PEArray.scala 200:17]
  wire [9:0] _GEN_330 = _T_24 ? 10'h0 : _GEN_127; // @[PEArray.scala 202:32 PEArray.scala 203:15]
  wire [2:0] _GEN_331 = _T_24 ? 3'h0 : state; // @[PEArray.scala 202:32 PEArray.scala 204:15 PEArray.scala 100:22]
  wire [9:0] _GEN_865 = {{4'd0}, GRU_out_width}; // @[PEArray.scala 220:19]
  wire [9:0] _GEN_0 = count % _GEN_865; // @[PEArray.scala 220:19]
  wire [5:0] _T_36 = _GEN_0[5:0]; // @[PEArray.scala 220:19]
  wire [5:0] _T_38 = GRU_out_width - 6'h1; // @[PEArray.scala 220:55]
  wire [5:0] _GEN_334 = _T_36 == _T_38 ? _L0Index_T_2 : 6'h0; // @[PEArray.scala 220:62 PEArray.scala 221:17 PEArray.scala 214:15]
  wire [5:0] _GEN_346 = _T_41 ? _GEN_334 : L0Index; // @[Conditional.scala 39:67 PEArray.scala 39:24]
  wire [9:0] _GEN_347 = _T_41 ? _GEN_330 : count; // @[Conditional.scala 39:67 PEArray.scala 101:22]
  wire [2:0] _GEN_348 = _T_41 ? _GEN_331 : state; // @[Conditional.scala 39:67 PEArray.scala 100:22]
  wire [5:0] _GEN_353 = _T_31 ? _GEN_334 : _GEN_346; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_354 = _T_31 ? _GEN_330 : _GEN_347; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_355 = _T_31 ? _GEN_331 : _GEN_348; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_356 = _T_22 ? _GEN_330 : _GEN_354; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_357 = _T_22 ? _GEN_329 : _GEN_353; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_458 = _T_22 ? _GEN_331 : _GEN_355; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_690 = _T_3 ? _GEN_118 : {{2'd0}, GRU_out_width}; // @[Conditional.scala 40:58 PEArray.scala 104:26]
  FP16MulAdder FP16MAC ( // @[PEArray.scala 72:23]
    .io_a(FP16MAC_io_a),
    .io_b(FP16MAC_io_b),
    .io_c(FP16MAC_io_c),
    .io_out(FP16MAC_io_out)
  );
  assign io_ToRightPE = mux3out_reg; // @[PEArray.scala 95:16]
  assign io_ToBelowPE = mux2out_reg; // @[PEArray.scala 94:16]
  assign FP16MAC_io_a = sel1 ? io_FromL1 : io_FromLeftPE; // @[PEArray.scala 50:14 PEArray.scala 50:23 PEArray.scala 51:24]
  assign FP16MAC_io_b = sel5 ? mux4out : _GEN_105; // @[PEArray.scala 77:13 PEArray.scala 78:18 PEArray.scala 81:18]
  assign FP16MAC_io_c = sel5 ? _GEN_105 : mux4out; // @[PEArray.scala 77:13 PEArray.scala 79:18 PEArray.scala 82:18]
  always @(posedge clock) begin
    if (reset) begin // @[PEArray.scala 39:24]
      L0Index <= 6'h0; // @[PEArray.scala 39:24]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h1; // @[PEArray.scala 159:15]
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h7; // @[PEArray.scala 181:15]
      end else begin
        L0Index <= _GEN_357;
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_0 <= _GEN_229;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_1 <= _GEN_230;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_2 <= _GEN_231;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_3 <= _GEN_232;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_4 <= _GEN_233;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_5 <= _GEN_234;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_6 <= _GEN_235;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_7 <= _GEN_236;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_8 <= _GEN_237;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_9 <= _GEN_238;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_10 <= _GEN_239;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_11 <= _GEN_240;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_12 <= _GEN_241;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_13 <= _GEN_242;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_14 <= _GEN_243;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_15 <= _GEN_244;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_16 <= _GEN_245;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_17 <= _GEN_246;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_18 <= _GEN_247;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_19 <= _GEN_248;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_20 <= _GEN_249;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_21 <= _GEN_250;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_22 <= _GEN_251;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_23 <= _GEN_252;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_24 <= _GEN_253;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_25 <= _GEN_254;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_26 <= _GEN_255;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_27 <= _GEN_256;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_28 <= _GEN_257;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_29 <= _GEN_258;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_30 <= _GEN_259;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_31 <= _GEN_260;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_32 <= _GEN_261;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_33 <= _GEN_262;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_34 <= _GEN_263;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_35 <= _GEN_264;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_36 <= _GEN_265;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_37 <= _GEN_266;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_38 <= _GEN_267;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_39 <= _GEN_268;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_40 <= _GEN_269;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_41 <= _GEN_270;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_42 <= _GEN_271;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_43 <= _GEN_272;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_44 <= _GEN_273;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_45 <= _GEN_274;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_46 <= _GEN_275;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_47 <= _GEN_276;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_48 <= _GEN_277;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_49 <= _GEN_278;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_50 <= _GEN_279;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_51 <= _GEN_280;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_52 <= _GEN_281;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_53 <= _GEN_282;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_54 <= _GEN_283;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_55 <= _GEN_284;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_56 <= _GEN_285;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_57 <= _GEN_286;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_58 <= _GEN_287;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_59 <= _GEN_288;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_60 <= _GEN_289;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_61 <= _GEN_290;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_62 <= _GEN_291;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_63 <= _GEN_292;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_64 <= _GEN_293;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_65 <= _GEN_294;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_66 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_67 <= _GEN_296;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_68 <= _GEN_297;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_69 <= _GEN_298;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_70 <= _GEN_299;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_71 <= _GEN_300;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_72 <= _GEN_301;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_73 <= _GEN_302;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_74 <= _GEN_303;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_75 <= _GEN_304;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_76 <= _GEN_305;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_77 <= _GEN_306;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_78 <= _GEN_307;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_79 <= _GEN_308;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_80 <= _GEN_309;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_81 <= _GEN_310;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_82 <= _GEN_311;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_83 <= _GEN_312;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_84 <= _GEN_313;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_85 <= _GEN_314;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_86 <= _GEN_315;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_87 <= _GEN_316;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_88 <= _GEN_317;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_89 <= _GEN_318;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_90 <= _GEN_319;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_91 <= _GEN_320;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_92 <= _GEN_321;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_93 <= _GEN_322;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_94 <= _GEN_323;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_95 <= _GEN_324;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_96 <= _GEN_325;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_97 <= _GEN_326;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_98 <= _GEN_327;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_99 <= _GEN_328;
          end
        end
      end
    end
    if (reset) begin // @[PEArray.scala 100:22]
      state <= 3'h0; // @[PEArray.scala 100:22]
    end else if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[7]) begin // @[PEArray.scala 116:57]
        state <= 3'h1;
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      if (count == 10'h33) begin // @[PEArray.scala 164:27]
        state <= 3'h0; // @[PEArray.scala 166:15]
      end
    end else if (_T_16) begin // @[Conditional.scala 39:67]
      state <= _GEN_126;
    end else begin
      state <= _GEN_458;
    end
    if (reset) begin // @[PEArray.scala 90:28]
      mux2out_reg <= 16'h0; // @[PEArray.scala 90:28]
    end else begin
      mux2out_reg <= MAC_out; // @[PEArray.scala 90:28]
    end
    if (reset) begin // @[PEArray.scala 91:28]
      mux3out_reg <= 16'h0; // @[PEArray.scala 91:28]
    end else if (sel3) begin // @[PEArray.scala 56:14]
      mux3out_reg <= MAC_out; // @[PEArray.scala 56:23]
    end else if (sel1) begin // @[PEArray.scala 50:14]
      mux3out_reg <= io_FromL1; // @[PEArray.scala 50:23]
    end else begin
      mux3out_reg <= io_FromLeftPE; // @[PEArray.scala 51:24]
    end
    if (reset) begin // @[PEArray.scala 101:22]
      count <= 10'h0; // @[PEArray.scala 101:22]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        if (count == 10'h33) begin // @[PEArray.scala 164:27]
          count <= 10'h0; // @[PEArray.scala 165:15]
        end else begin
          count <= _GEN_120;
        end
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        count <= _GEN_125;
      end else begin
        count <= _GEN_356;
      end
    end
    GRU_out_width <= _GEN_690[5:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  L0Index = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  L0Memory_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  L0Memory_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  L0Memory_2 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  L0Memory_3 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  L0Memory_4 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  L0Memory_5 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  L0Memory_6 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  L0Memory_7 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  L0Memory_8 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  L0Memory_9 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  L0Memory_10 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  L0Memory_11 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  L0Memory_12 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  L0Memory_13 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  L0Memory_14 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  L0Memory_15 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  L0Memory_16 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  L0Memory_17 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  L0Memory_18 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  L0Memory_19 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  L0Memory_20 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  L0Memory_21 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  L0Memory_22 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  L0Memory_23 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  L0Memory_24 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  L0Memory_25 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  L0Memory_26 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  L0Memory_27 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  L0Memory_28 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  L0Memory_29 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  L0Memory_30 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  L0Memory_31 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  L0Memory_32 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  L0Memory_33 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  L0Memory_34 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  L0Memory_35 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  L0Memory_36 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  L0Memory_37 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  L0Memory_38 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  L0Memory_39 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  L0Memory_40 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  L0Memory_41 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  L0Memory_42 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  L0Memory_43 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  L0Memory_44 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  L0Memory_45 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  L0Memory_46 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  L0Memory_47 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  L0Memory_48 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  L0Memory_49 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  L0Memory_50 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  L0Memory_51 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  L0Memory_52 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  L0Memory_53 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  L0Memory_54 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  L0Memory_55 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  L0Memory_56 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  L0Memory_57 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  L0Memory_58 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  L0Memory_59 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  L0Memory_60 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  L0Memory_61 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  L0Memory_62 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  L0Memory_63 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  L0Memory_64 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  L0Memory_65 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  L0Memory_66 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  L0Memory_67 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  L0Memory_68 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  L0Memory_69 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  L0Memory_70 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  L0Memory_71 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  L0Memory_72 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  L0Memory_73 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  L0Memory_74 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  L0Memory_75 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  L0Memory_76 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  L0Memory_77 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  L0Memory_78 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  L0Memory_79 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  L0Memory_80 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  L0Memory_81 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  L0Memory_82 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  L0Memory_83 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  L0Memory_84 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  L0Memory_85 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  L0Memory_86 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  L0Memory_87 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  L0Memory_88 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  L0Memory_89 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  L0Memory_90 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  L0Memory_91 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  L0Memory_92 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  L0Memory_93 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  L0Memory_94 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  L0Memory_95 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  L0Memory_96 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  L0Memory_97 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  L0Memory_98 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  L0Memory_99 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  state = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  mux2out_reg = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  mux3out_reg = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  count = _RAND_104[9:0];
  _RAND_105 = {1{`RANDOM}};
  GRU_out_width = _RAND_105[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PE_14(
  input         clock,
  input         reset,
  input  [15:0] io_FromAbovePE,
  input  [15:0] io_FromLeftPE,
  input  [15:0] io_FromL1,
  input  [2:0]  io_control_signal_control,
  input  [9:0]  io_control_signal_count,
  input  [5:0]  io_control_signal_L0index,
  input  [11:0] io_control_signal_mask,
  input  [7:0]  io_control_signal_gru_out_width,
  output [15:0] io_ToRightPE,
  output [15:0] io_ToBelowPE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] FP16MAC_io_a; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_b; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_c; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_out; // @[PEArray.scala 72:23]
  reg [5:0] L0Index; // @[PEArray.scala 39:24]
  reg [15:0] L0Memory_0; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_1; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_2; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_3; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_4; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_5; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_6; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_7; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_8; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_9; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_10; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_11; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_12; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_13; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_14; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_15; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_16; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_17; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_18; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_19; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_20; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_21; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_22; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_23; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_24; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_25; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_26; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_27; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_28; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_29; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_30; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_31; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_32; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_33; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_34; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_35; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_36; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_37; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_38; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_39; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_40; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_41; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_42; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_43; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_44; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_45; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_46; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_47; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_48; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_49; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_50; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_51; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_52; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_53; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_54; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_55; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_56; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_57; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_58; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_59; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_60; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_61; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_62; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_63; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_64; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_65; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_66; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_67; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_68; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_69; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_70; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_71; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_72; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_73; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_74; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_75; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_76; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_77; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_78; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_79; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_80; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_81; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_82; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_83; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_84; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_85; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_86; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_87; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_88; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_89; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_90; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_91; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_92; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_93; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_94; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_95; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_96; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_97; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_98; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_99; // @[PEArray.scala 40:21]
  reg [2:0] state; // @[PEArray.scala 100:22]
  wire  _T_3 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_12 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_16 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_22 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_31 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_41 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_342 = _T_41 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 231:12 PEArray.scala 32:8]
  wire  _GEN_349 = _T_31 ? 1'h0 : _GEN_342; // @[Conditional.scala 39:67 PEArray.scala 208:12]
  wire  _GEN_459 = _T_22 | _GEN_349; // @[Conditional.scala 39:67 PEArray.scala 32:8]
  wire  _GEN_463 = _T_16 ? 1'h0 : _GEN_459; // @[Conditional.scala 39:67]
  wire  _GEN_572 = _T_12 | _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 149:12]
  wire  sel1 = _T_3 | _GEN_572; // @[Conditional.scala 40:58 PEArray.scala 108:12]
  wire [15:0] MAC_out = FP16MAC_io_out; // @[PEArray.scala 47:21 PEArray.scala 85:11]
  wire  _GEN_465 = _T_16 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 177:12]
  wire  _GEN_580 = _T_12 | _GEN_465; // @[Conditional.scala 39:67 PEArray.scala 34:8]
  wire  sel3 = _T_3 | _GEN_580; // @[Conditional.scala 40:58 PEArray.scala 110:12]
  wire [1:0] _GEN_344 = _T_41 ? 2'h2 : 2'h0; // @[Conditional.scala 39:67 PEArray.scala 233:12 PEArray.scala 35:8]
  wire [1:0] _GEN_351 = _T_31 ? 2'h2 : _GEN_344; // @[Conditional.scala 39:67 PEArray.scala 210:12]
  wire [1:0] _GEN_461 = _T_22 ? 2'h0 : _GEN_351; // @[Conditional.scala 39:67 PEArray.scala 35:8]
  wire [1:0] _GEN_466 = _T_16 ? 2'h0 : _GEN_461; // @[Conditional.scala 39:67 PEArray.scala 178:12]
  wire [1:0] _GEN_574 = _T_12 ? 2'h1 : _GEN_466; // @[Conditional.scala 39:67]
  wire [1:0] sel4 = _T_3 ? 2'h0 : _GEN_574; // @[Conditional.scala 40:58 PEArray.scala 111:12]
  wire [15:0] _GEN_3 = sel4 == 2'h2 ? io_FromL1 : 16'h0; // @[PEArray.scala 65:28 PEArray.scala 66:15 PEArray.scala 69:15]
  wire [15:0] _GEN_4 = sel4 == 2'h1 ? io_FromAbovePE : _GEN_3; // @[PEArray.scala 62:28 PEArray.scala 63:15]
  wire [15:0] mux4out = sel4 == 2'h0 ? 16'h0 : _GEN_4; // @[PEArray.scala 59:22 PEArray.scala 60:13]
  wire [15:0] _GEN_7 = 6'h1 == L0Index ? L0Memory_1 : L0Memory_0; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_8 = 6'h2 == L0Index ? L0Memory_2 : _GEN_7; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_9 = 6'h3 == L0Index ? L0Memory_3 : _GEN_8; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_10 = 6'h4 == L0Index ? L0Memory_4 : _GEN_9; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_11 = 6'h5 == L0Index ? L0Memory_5 : _GEN_10; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_12 = 6'h6 == L0Index ? L0Memory_6 : _GEN_11; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_13 = 6'h7 == L0Index ? L0Memory_7 : _GEN_12; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_14 = 6'h8 == L0Index ? L0Memory_8 : _GEN_13; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_15 = 6'h9 == L0Index ? L0Memory_9 : _GEN_14; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_16 = 6'ha == L0Index ? L0Memory_10 : _GEN_15; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_17 = 6'hb == L0Index ? L0Memory_11 : _GEN_16; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_18 = 6'hc == L0Index ? L0Memory_12 : _GEN_17; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_19 = 6'hd == L0Index ? L0Memory_13 : _GEN_18; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_20 = 6'he == L0Index ? L0Memory_14 : _GEN_19; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_21 = 6'hf == L0Index ? L0Memory_15 : _GEN_20; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_22 = 6'h10 == L0Index ? L0Memory_16 : _GEN_21; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_23 = 6'h11 == L0Index ? L0Memory_17 : _GEN_22; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_24 = 6'h12 == L0Index ? L0Memory_18 : _GEN_23; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_25 = 6'h13 == L0Index ? L0Memory_19 : _GEN_24; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_26 = 6'h14 == L0Index ? L0Memory_20 : _GEN_25; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_27 = 6'h15 == L0Index ? L0Memory_21 : _GEN_26; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_28 = 6'h16 == L0Index ? L0Memory_22 : _GEN_27; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_29 = 6'h17 == L0Index ? L0Memory_23 : _GEN_28; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_30 = 6'h18 == L0Index ? L0Memory_24 : _GEN_29; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_31 = 6'h19 == L0Index ? L0Memory_25 : _GEN_30; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_32 = 6'h1a == L0Index ? L0Memory_26 : _GEN_31; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_33 = 6'h1b == L0Index ? L0Memory_27 : _GEN_32; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_34 = 6'h1c == L0Index ? L0Memory_28 : _GEN_33; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_35 = 6'h1d == L0Index ? L0Memory_29 : _GEN_34; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_36 = 6'h1e == L0Index ? L0Memory_30 : _GEN_35; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_37 = 6'h1f == L0Index ? L0Memory_31 : _GEN_36; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_38 = 6'h20 == L0Index ? L0Memory_32 : _GEN_37; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_39 = 6'h21 == L0Index ? L0Memory_33 : _GEN_38; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_40 = 6'h22 == L0Index ? L0Memory_34 : _GEN_39; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_41 = 6'h23 == L0Index ? L0Memory_35 : _GEN_40; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_42 = 6'h24 == L0Index ? L0Memory_36 : _GEN_41; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_43 = 6'h25 == L0Index ? L0Memory_37 : _GEN_42; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_44 = 6'h26 == L0Index ? L0Memory_38 : _GEN_43; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_45 = 6'h27 == L0Index ? L0Memory_39 : _GEN_44; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_46 = 6'h28 == L0Index ? L0Memory_40 : _GEN_45; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_47 = 6'h29 == L0Index ? L0Memory_41 : _GEN_46; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_48 = 6'h2a == L0Index ? L0Memory_42 : _GEN_47; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_49 = 6'h2b == L0Index ? L0Memory_43 : _GEN_48; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_50 = 6'h2c == L0Index ? L0Memory_44 : _GEN_49; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_51 = 6'h2d == L0Index ? L0Memory_45 : _GEN_50; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_52 = 6'h2e == L0Index ? L0Memory_46 : _GEN_51; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_53 = 6'h2f == L0Index ? L0Memory_47 : _GEN_52; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_54 = 6'h30 == L0Index ? L0Memory_48 : _GEN_53; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_55 = 6'h31 == L0Index ? L0Memory_49 : _GEN_54; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_56 = 6'h32 == L0Index ? L0Memory_50 : _GEN_55; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_57 = 6'h33 == L0Index ? L0Memory_51 : _GEN_56; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_58 = 6'h34 == L0Index ? L0Memory_52 : _GEN_57; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_59 = 6'h35 == L0Index ? L0Memory_53 : _GEN_58; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_60 = 6'h36 == L0Index ? L0Memory_54 : _GEN_59; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_61 = 6'h37 == L0Index ? L0Memory_55 : _GEN_60; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_62 = 6'h38 == L0Index ? L0Memory_56 : _GEN_61; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_63 = 6'h39 == L0Index ? L0Memory_57 : _GEN_62; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_64 = 6'h3a == L0Index ? L0Memory_58 : _GEN_63; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_65 = 6'h3b == L0Index ? L0Memory_59 : _GEN_64; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_66 = 6'h3c == L0Index ? L0Memory_60 : _GEN_65; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_67 = 6'h3d == L0Index ? L0Memory_61 : _GEN_66; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_68 = 6'h3e == L0Index ? L0Memory_62 : _GEN_67; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_69 = 6'h3f == L0Index ? L0Memory_63 : _GEN_68; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [6:0] _GEN_793 = {{1'd0}, L0Index}; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_70 = 7'h40 == _GEN_793 ? L0Memory_64 : _GEN_69; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_71 = 7'h41 == _GEN_793 ? L0Memory_65 : _GEN_70; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_72 = 7'h42 == _GEN_793 ? L0Memory_66 : _GEN_71; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_73 = 7'h43 == _GEN_793 ? L0Memory_67 : _GEN_72; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_74 = 7'h44 == _GEN_793 ? L0Memory_68 : _GEN_73; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_75 = 7'h45 == _GEN_793 ? L0Memory_69 : _GEN_74; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_76 = 7'h46 == _GEN_793 ? L0Memory_70 : _GEN_75; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_77 = 7'h47 == _GEN_793 ? L0Memory_71 : _GEN_76; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_78 = 7'h48 == _GEN_793 ? L0Memory_72 : _GEN_77; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_79 = 7'h49 == _GEN_793 ? L0Memory_73 : _GEN_78; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_80 = 7'h4a == _GEN_793 ? L0Memory_74 : _GEN_79; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_81 = 7'h4b == _GEN_793 ? L0Memory_75 : _GEN_80; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_82 = 7'h4c == _GEN_793 ? L0Memory_76 : _GEN_81; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_83 = 7'h4d == _GEN_793 ? L0Memory_77 : _GEN_82; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_84 = 7'h4e == _GEN_793 ? L0Memory_78 : _GEN_83; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_85 = 7'h4f == _GEN_793 ? L0Memory_79 : _GEN_84; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_86 = 7'h50 == _GEN_793 ? L0Memory_80 : _GEN_85; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_87 = 7'h51 == _GEN_793 ? L0Memory_81 : _GEN_86; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_88 = 7'h52 == _GEN_793 ? L0Memory_82 : _GEN_87; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_89 = 7'h53 == _GEN_793 ? L0Memory_83 : _GEN_88; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_90 = 7'h54 == _GEN_793 ? L0Memory_84 : _GEN_89; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_91 = 7'h55 == _GEN_793 ? L0Memory_85 : _GEN_90; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_92 = 7'h56 == _GEN_793 ? L0Memory_86 : _GEN_91; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_93 = 7'h57 == _GEN_793 ? L0Memory_87 : _GEN_92; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_94 = 7'h58 == _GEN_793 ? L0Memory_88 : _GEN_93; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_95 = 7'h59 == _GEN_793 ? L0Memory_89 : _GEN_94; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_96 = 7'h5a == _GEN_793 ? L0Memory_90 : _GEN_95; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_97 = 7'h5b == _GEN_793 ? L0Memory_91 : _GEN_96; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_98 = 7'h5c == _GEN_793 ? L0Memory_92 : _GEN_97; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_99 = 7'h5d == _GEN_793 ? L0Memory_93 : _GEN_98; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_100 = 7'h5e == _GEN_793 ? L0Memory_94 : _GEN_99; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_101 = 7'h5f == _GEN_793 ? L0Memory_95 : _GEN_100; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_102 = 7'h60 == _GEN_793 ? L0Memory_96 : _GEN_101; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_103 = 7'h61 == _GEN_793 ? L0Memory_97 : _GEN_102; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_104 = 7'h62 == _GEN_793 ? L0Memory_98 : _GEN_103; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_105 = 7'h63 == _GEN_793 ? L0Memory_99 : _GEN_104; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire  _GEN_575 = _T_12 ? 1'h0 : _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 157:12]
  wire  sel5 = _T_3 ? 1'h0 : _GEN_575; // @[Conditional.scala 40:58 PEArray.scala 112:12]
  reg [15:0] mux2out_reg; // @[PEArray.scala 90:28]
  reg [15:0] mux3out_reg; // @[PEArray.scala 91:28]
  reg [9:0] count; // @[PEArray.scala 101:22]
  reg [9:0] count_max; // @[PEArray.scala 102:22]
  reg [5:0] L0index_begin; // @[PEArray.scala 103:26]
  reg [5:0] GRU_out_width; // @[PEArray.scala 104:26]
  wire  _T_6 = 3'h0 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_7 = 3'h1 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_8 = 3'h2 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_9 = 3'h3 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_10 = 3'h4 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_11 = 3'h5 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_109 = _T_11 ? 3'h5 : state; // @[Conditional.scala 39:67 PEArray.scala 140:19 PEArray.scala 100:22]
  wire [2:0] _GEN_110 = _T_10 ? 3'h4 : _GEN_109; // @[Conditional.scala 39:67 PEArray.scala 136:19]
  wire [2:0] _GEN_111 = _T_9 ? 3'h3 : _GEN_110; // @[Conditional.scala 39:67 PEArray.scala 132:19]
  wire [2:0] _GEN_112 = _T_8 ? 3'h2 : _GEN_111; // @[Conditional.scala 39:67 PEArray.scala 128:19]
  wire [2:0] _GEN_113 = _T_7 ? 3'h1 : _GEN_112; // @[Conditional.scala 39:67 PEArray.scala 124:19]
  wire [7:0] _GEN_118 = io_control_signal_mask[7] ? io_control_signal_gru_out_width : {{2'd0}, GRU_out_width}; // @[PEArray.scala 116:57 PEArray.scala 145:23 PEArray.scala 104:26]
  wire [9:0] _count_T_1 = count + 10'h1; // @[PEArray.scala 162:24]
  wire [9:0] _GEN_120 = count != 10'h33 ? _count_T_1 : count; // @[PEArray.scala 161:27 PEArray.scala 162:15 PEArray.scala 101:22]
  wire [9:0] _GEN_124 = count != 10'h188 ? _count_T_1 : count; // @[PEArray.scala 183:28 PEArray.scala 184:15 PEArray.scala 101:22]
  wire [9:0] _GEN_125 = count == 10'h188 ? 10'h0 : _GEN_124; // @[PEArray.scala 186:28 PEArray.scala 187:15]
  wire [2:0] _GEN_126 = count == 10'h188 ? 3'h0 : state; // @[PEArray.scala 186:28 PEArray.scala 188:15 PEArray.scala 100:22]
  wire [9:0] _GEN_127 = count != count_max ? _count_T_1 : count; // @[PEArray.scala 192:32 PEArray.scala 193:15 PEArray.scala 101:22]
  wire [5:0] _GEN_128 = count == 10'h0 ? L0index_begin : L0Index; // @[PEArray.scala 195:26 PEArray.scala 196:17 PEArray.scala 39:24]
  wire [9:0] _T_27 = count_max - 10'h1; // @[PEArray.scala 198:51]
  wire [15:0] _GEN_129 = 6'h0 == L0Index ? io_FromL1 : L0Memory_0; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_130 = 6'h1 == L0Index ? io_FromL1 : L0Memory_1; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_131 = 6'h2 == L0Index ? io_FromL1 : L0Memory_2; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_132 = 6'h3 == L0Index ? io_FromL1 : L0Memory_3; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_133 = 6'h4 == L0Index ? io_FromL1 : L0Memory_4; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_134 = 6'h5 == L0Index ? io_FromL1 : L0Memory_5; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_135 = 6'h6 == L0Index ? io_FromL1 : L0Memory_6; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_136 = 6'h7 == L0Index ? io_FromL1 : L0Memory_7; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_137 = 6'h8 == L0Index ? io_FromL1 : L0Memory_8; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_138 = 6'h9 == L0Index ? io_FromL1 : L0Memory_9; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_139 = 6'ha == L0Index ? io_FromL1 : L0Memory_10; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_140 = 6'hb == L0Index ? io_FromL1 : L0Memory_11; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_141 = 6'hc == L0Index ? io_FromL1 : L0Memory_12; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_142 = 6'hd == L0Index ? io_FromL1 : L0Memory_13; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_143 = 6'he == L0Index ? io_FromL1 : L0Memory_14; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_144 = 6'hf == L0Index ? io_FromL1 : L0Memory_15; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_145 = 6'h10 == L0Index ? io_FromL1 : L0Memory_16; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_146 = 6'h11 == L0Index ? io_FromL1 : L0Memory_17; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_147 = 6'h12 == L0Index ? io_FromL1 : L0Memory_18; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_148 = 6'h13 == L0Index ? io_FromL1 : L0Memory_19; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_149 = 6'h14 == L0Index ? io_FromL1 : L0Memory_20; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_150 = 6'h15 == L0Index ? io_FromL1 : L0Memory_21; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_151 = 6'h16 == L0Index ? io_FromL1 : L0Memory_22; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_152 = 6'h17 == L0Index ? io_FromL1 : L0Memory_23; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_153 = 6'h18 == L0Index ? io_FromL1 : L0Memory_24; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_154 = 6'h19 == L0Index ? io_FromL1 : L0Memory_25; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_155 = 6'h1a == L0Index ? io_FromL1 : L0Memory_26; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_156 = 6'h1b == L0Index ? io_FromL1 : L0Memory_27; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_157 = 6'h1c == L0Index ? io_FromL1 : L0Memory_28; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_158 = 6'h1d == L0Index ? io_FromL1 : L0Memory_29; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_159 = 6'h1e == L0Index ? io_FromL1 : L0Memory_30; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_160 = 6'h1f == L0Index ? io_FromL1 : L0Memory_31; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_161 = 6'h20 == L0Index ? io_FromL1 : L0Memory_32; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_162 = 6'h21 == L0Index ? io_FromL1 : L0Memory_33; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_163 = 6'h22 == L0Index ? io_FromL1 : L0Memory_34; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_164 = 6'h23 == L0Index ? io_FromL1 : L0Memory_35; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_165 = 6'h24 == L0Index ? io_FromL1 : L0Memory_36; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_166 = 6'h25 == L0Index ? io_FromL1 : L0Memory_37; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_167 = 6'h26 == L0Index ? io_FromL1 : L0Memory_38; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_168 = 6'h27 == L0Index ? io_FromL1 : L0Memory_39; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_169 = 6'h28 == L0Index ? io_FromL1 : L0Memory_40; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_170 = 6'h29 == L0Index ? io_FromL1 : L0Memory_41; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_171 = 6'h2a == L0Index ? io_FromL1 : L0Memory_42; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_172 = 6'h2b == L0Index ? io_FromL1 : L0Memory_43; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_173 = 6'h2c == L0Index ? io_FromL1 : L0Memory_44; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_174 = 6'h2d == L0Index ? io_FromL1 : L0Memory_45; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_175 = 6'h2e == L0Index ? io_FromL1 : L0Memory_46; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_176 = 6'h2f == L0Index ? io_FromL1 : L0Memory_47; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_177 = 6'h30 == L0Index ? io_FromL1 : L0Memory_48; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_178 = 6'h31 == L0Index ? io_FromL1 : L0Memory_49; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_179 = 6'h32 == L0Index ? io_FromL1 : L0Memory_50; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_180 = 6'h33 == L0Index ? io_FromL1 : L0Memory_51; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_181 = 6'h34 == L0Index ? io_FromL1 : L0Memory_52; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_182 = 6'h35 == L0Index ? io_FromL1 : L0Memory_53; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_183 = 6'h36 == L0Index ? io_FromL1 : L0Memory_54; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_184 = 6'h37 == L0Index ? io_FromL1 : L0Memory_55; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_185 = 6'h38 == L0Index ? io_FromL1 : L0Memory_56; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_186 = 6'h39 == L0Index ? io_FromL1 : L0Memory_57; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_187 = 6'h3a == L0Index ? io_FromL1 : L0Memory_58; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_188 = 6'h3b == L0Index ? io_FromL1 : L0Memory_59; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_189 = 6'h3c == L0Index ? io_FromL1 : L0Memory_60; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_190 = 6'h3d == L0Index ? io_FromL1 : L0Memory_61; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_191 = 6'h3e == L0Index ? io_FromL1 : L0Memory_62; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_192 = 6'h3f == L0Index ? io_FromL1 : L0Memory_63; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_193 = 7'h40 == _GEN_793 ? io_FromL1 : L0Memory_64; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_194 = 7'h41 == _GEN_793 ? io_FromL1 : L0Memory_65; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_195 = 7'h42 == _GEN_793 ? io_FromL1 : L0Memory_66; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_196 = 7'h43 == _GEN_793 ? io_FromL1 : L0Memory_67; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_197 = 7'h44 == _GEN_793 ? io_FromL1 : L0Memory_68; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_198 = 7'h45 == _GEN_793 ? io_FromL1 : L0Memory_69; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_199 = 7'h46 == _GEN_793 ? io_FromL1 : L0Memory_70; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_200 = 7'h47 == _GEN_793 ? io_FromL1 : L0Memory_71; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_201 = 7'h48 == _GEN_793 ? io_FromL1 : L0Memory_72; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_202 = 7'h49 == _GEN_793 ? io_FromL1 : L0Memory_73; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_203 = 7'h4a == _GEN_793 ? io_FromL1 : L0Memory_74; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_204 = 7'h4b == _GEN_793 ? io_FromL1 : L0Memory_75; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_205 = 7'h4c == _GEN_793 ? io_FromL1 : L0Memory_76; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_206 = 7'h4d == _GEN_793 ? io_FromL1 : L0Memory_77; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_207 = 7'h4e == _GEN_793 ? io_FromL1 : L0Memory_78; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_208 = 7'h4f == _GEN_793 ? io_FromL1 : L0Memory_79; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_209 = 7'h50 == _GEN_793 ? io_FromL1 : L0Memory_80; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_210 = 7'h51 == _GEN_793 ? io_FromL1 : L0Memory_81; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_211 = 7'h52 == _GEN_793 ? io_FromL1 : L0Memory_82; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_212 = 7'h53 == _GEN_793 ? io_FromL1 : L0Memory_83; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_213 = 7'h54 == _GEN_793 ? io_FromL1 : L0Memory_84; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_214 = 7'h55 == _GEN_793 ? io_FromL1 : L0Memory_85; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_215 = 7'h56 == _GEN_793 ? io_FromL1 : L0Memory_86; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_216 = 7'h57 == _GEN_793 ? io_FromL1 : L0Memory_87; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_217 = 7'h58 == _GEN_793 ? io_FromL1 : L0Memory_88; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_218 = 7'h59 == _GEN_793 ? io_FromL1 : L0Memory_89; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_219 = 7'h5a == _GEN_793 ? io_FromL1 : L0Memory_90; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_220 = 7'h5b == _GEN_793 ? io_FromL1 : L0Memory_91; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_221 = 7'h5c == _GEN_793 ? io_FromL1 : L0Memory_92; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_222 = 7'h5d == _GEN_793 ? io_FromL1 : L0Memory_93; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_223 = 7'h5e == _GEN_793 ? io_FromL1 : L0Memory_94; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_224 = 7'h5f == _GEN_793 ? io_FromL1 : L0Memory_95; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_225 = 7'h60 == _GEN_793 ? io_FromL1 : L0Memory_96; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_226 = 7'h61 == _GEN_793 ? io_FromL1 : L0Memory_97; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_227 = 7'h62 == _GEN_793 ? io_FromL1 : L0Memory_98; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_228 = 7'h63 == _GEN_793 ? io_FromL1 : L0Memory_99; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [5:0] _L0Index_T_2 = L0Index + 6'h1; // @[PEArray.scala 200:28]
  wire [15:0] _GEN_229 = count >= 10'h1 & count <= _T_27 ? _GEN_129 : L0Memory_0; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_230 = count >= 10'h1 & count <= _T_27 ? _GEN_130 : L0Memory_1; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_231 = count >= 10'h1 & count <= _T_27 ? _GEN_131 : L0Memory_2; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_232 = count >= 10'h1 & count <= _T_27 ? _GEN_132 : L0Memory_3; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_233 = count >= 10'h1 & count <= _T_27 ? _GEN_133 : L0Memory_4; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_234 = count >= 10'h1 & count <= _T_27 ? _GEN_134 : L0Memory_5; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_235 = count >= 10'h1 & count <= _T_27 ? _GEN_135 : L0Memory_6; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_236 = count >= 10'h1 & count <= _T_27 ? _GEN_136 : L0Memory_7; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_237 = count >= 10'h1 & count <= _T_27 ? _GEN_137 : L0Memory_8; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_238 = count >= 10'h1 & count <= _T_27 ? _GEN_138 : L0Memory_9; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_239 = count >= 10'h1 & count <= _T_27 ? _GEN_139 : L0Memory_10; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_240 = count >= 10'h1 & count <= _T_27 ? _GEN_140 : L0Memory_11; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_241 = count >= 10'h1 & count <= _T_27 ? _GEN_141 : L0Memory_12; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_242 = count >= 10'h1 & count <= _T_27 ? _GEN_142 : L0Memory_13; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_243 = count >= 10'h1 & count <= _T_27 ? _GEN_143 : L0Memory_14; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_244 = count >= 10'h1 & count <= _T_27 ? _GEN_144 : L0Memory_15; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_245 = count >= 10'h1 & count <= _T_27 ? _GEN_145 : L0Memory_16; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_246 = count >= 10'h1 & count <= _T_27 ? _GEN_146 : L0Memory_17; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_247 = count >= 10'h1 & count <= _T_27 ? _GEN_147 : L0Memory_18; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_248 = count >= 10'h1 & count <= _T_27 ? _GEN_148 : L0Memory_19; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_249 = count >= 10'h1 & count <= _T_27 ? _GEN_149 : L0Memory_20; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_250 = count >= 10'h1 & count <= _T_27 ? _GEN_150 : L0Memory_21; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_251 = count >= 10'h1 & count <= _T_27 ? _GEN_151 : L0Memory_22; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_252 = count >= 10'h1 & count <= _T_27 ? _GEN_152 : L0Memory_23; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_253 = count >= 10'h1 & count <= _T_27 ? _GEN_153 : L0Memory_24; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_254 = count >= 10'h1 & count <= _T_27 ? _GEN_154 : L0Memory_25; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_255 = count >= 10'h1 & count <= _T_27 ? _GEN_155 : L0Memory_26; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_256 = count >= 10'h1 & count <= _T_27 ? _GEN_156 : L0Memory_27; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_257 = count >= 10'h1 & count <= _T_27 ? _GEN_157 : L0Memory_28; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_258 = count >= 10'h1 & count <= _T_27 ? _GEN_158 : L0Memory_29; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_259 = count >= 10'h1 & count <= _T_27 ? _GEN_159 : L0Memory_30; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_260 = count >= 10'h1 & count <= _T_27 ? _GEN_160 : L0Memory_31; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_261 = count >= 10'h1 & count <= _T_27 ? _GEN_161 : L0Memory_32; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_262 = count >= 10'h1 & count <= _T_27 ? _GEN_162 : L0Memory_33; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_263 = count >= 10'h1 & count <= _T_27 ? _GEN_163 : L0Memory_34; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_264 = count >= 10'h1 & count <= _T_27 ? _GEN_164 : L0Memory_35; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_265 = count >= 10'h1 & count <= _T_27 ? _GEN_165 : L0Memory_36; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_266 = count >= 10'h1 & count <= _T_27 ? _GEN_166 : L0Memory_37; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_267 = count >= 10'h1 & count <= _T_27 ? _GEN_167 : L0Memory_38; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_268 = count >= 10'h1 & count <= _T_27 ? _GEN_168 : L0Memory_39; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_269 = count >= 10'h1 & count <= _T_27 ? _GEN_169 : L0Memory_40; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_270 = count >= 10'h1 & count <= _T_27 ? _GEN_170 : L0Memory_41; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_271 = count >= 10'h1 & count <= _T_27 ? _GEN_171 : L0Memory_42; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_272 = count >= 10'h1 & count <= _T_27 ? _GEN_172 : L0Memory_43; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_273 = count >= 10'h1 & count <= _T_27 ? _GEN_173 : L0Memory_44; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_274 = count >= 10'h1 & count <= _T_27 ? _GEN_174 : L0Memory_45; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_275 = count >= 10'h1 & count <= _T_27 ? _GEN_175 : L0Memory_46; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_276 = count >= 10'h1 & count <= _T_27 ? _GEN_176 : L0Memory_47; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_277 = count >= 10'h1 & count <= _T_27 ? _GEN_177 : L0Memory_48; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_278 = count >= 10'h1 & count <= _T_27 ? _GEN_178 : L0Memory_49; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_279 = count >= 10'h1 & count <= _T_27 ? _GEN_179 : L0Memory_50; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_280 = count >= 10'h1 & count <= _T_27 ? _GEN_180 : L0Memory_51; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_281 = count >= 10'h1 & count <= _T_27 ? _GEN_181 : L0Memory_52; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_282 = count >= 10'h1 & count <= _T_27 ? _GEN_182 : L0Memory_53; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_283 = count >= 10'h1 & count <= _T_27 ? _GEN_183 : L0Memory_54; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_284 = count >= 10'h1 & count <= _T_27 ? _GEN_184 : L0Memory_55; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_285 = count >= 10'h1 & count <= _T_27 ? _GEN_185 : L0Memory_56; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_286 = count >= 10'h1 & count <= _T_27 ? _GEN_186 : L0Memory_57; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_287 = count >= 10'h1 & count <= _T_27 ? _GEN_187 : L0Memory_58; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_288 = count >= 10'h1 & count <= _T_27 ? _GEN_188 : L0Memory_59; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_289 = count >= 10'h1 & count <= _T_27 ? _GEN_189 : L0Memory_60; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_290 = count >= 10'h1 & count <= _T_27 ? _GEN_190 : L0Memory_61; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_291 = count >= 10'h1 & count <= _T_27 ? _GEN_191 : L0Memory_62; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_292 = count >= 10'h1 & count <= _T_27 ? _GEN_192 : L0Memory_63; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_293 = count >= 10'h1 & count <= _T_27 ? _GEN_193 : L0Memory_64; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_294 = count >= 10'h1 & count <= _T_27 ? _GEN_194 : L0Memory_65; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_295 = count >= 10'h1 & count <= _T_27 ? _GEN_195 : L0Memory_66; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_296 = count >= 10'h1 & count <= _T_27 ? _GEN_196 : L0Memory_67; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_297 = count >= 10'h1 & count <= _T_27 ? _GEN_197 : L0Memory_68; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_298 = count >= 10'h1 & count <= _T_27 ? _GEN_198 : L0Memory_69; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_299 = count >= 10'h1 & count <= _T_27 ? _GEN_199 : L0Memory_70; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_300 = count >= 10'h1 & count <= _T_27 ? _GEN_200 : L0Memory_71; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_301 = count >= 10'h1 & count <= _T_27 ? _GEN_201 : L0Memory_72; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_302 = count >= 10'h1 & count <= _T_27 ? _GEN_202 : L0Memory_73; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_303 = count >= 10'h1 & count <= _T_27 ? _GEN_203 : L0Memory_74; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_304 = count >= 10'h1 & count <= _T_27 ? _GEN_204 : L0Memory_75; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_305 = count >= 10'h1 & count <= _T_27 ? _GEN_205 : L0Memory_76; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_306 = count >= 10'h1 & count <= _T_27 ? _GEN_206 : L0Memory_77; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_307 = count >= 10'h1 & count <= _T_27 ? _GEN_207 : L0Memory_78; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_308 = count >= 10'h1 & count <= _T_27 ? _GEN_208 : L0Memory_79; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_309 = count >= 10'h1 & count <= _T_27 ? _GEN_209 : L0Memory_80; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_310 = count >= 10'h1 & count <= _T_27 ? _GEN_210 : L0Memory_81; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_311 = count >= 10'h1 & count <= _T_27 ? _GEN_211 : L0Memory_82; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_312 = count >= 10'h1 & count <= _T_27 ? _GEN_212 : L0Memory_83; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_313 = count >= 10'h1 & count <= _T_27 ? _GEN_213 : L0Memory_84; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_314 = count >= 10'h1 & count <= _T_27 ? _GEN_214 : L0Memory_85; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_315 = count >= 10'h1 & count <= _T_27 ? _GEN_215 : L0Memory_86; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_316 = count >= 10'h1 & count <= _T_27 ? _GEN_216 : L0Memory_87; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_317 = count >= 10'h1 & count <= _T_27 ? _GEN_217 : L0Memory_88; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_318 = count >= 10'h1 & count <= _T_27 ? _GEN_218 : L0Memory_89; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_319 = count >= 10'h1 & count <= _T_27 ? _GEN_219 : L0Memory_90; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_320 = count >= 10'h1 & count <= _T_27 ? _GEN_220 : L0Memory_91; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_321 = count >= 10'h1 & count <= _T_27 ? _GEN_221 : L0Memory_92; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_322 = count >= 10'h1 & count <= _T_27 ? _GEN_222 : L0Memory_93; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_323 = count >= 10'h1 & count <= _T_27 ? _GEN_223 : L0Memory_94; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_324 = count >= 10'h1 & count <= _T_27 ? _GEN_224 : L0Memory_95; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_325 = count >= 10'h1 & count <= _T_27 ? _GEN_225 : L0Memory_96; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_326 = count >= 10'h1 & count <= _T_27 ? _GEN_226 : L0Memory_97; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_327 = count >= 10'h1 & count <= _T_27 ? _GEN_227 : L0Memory_98; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_328 = count >= 10'h1 & count <= _T_27 ? _GEN_228 : L0Memory_99; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [5:0] _GEN_329 = count >= 10'h1 & count <= _T_27 ? _L0Index_T_2 : _GEN_128; // @[PEArray.scala 198:59 PEArray.scala 200:17]
  wire [9:0] _GEN_330 = count == count_max ? 10'h0 : _GEN_127; // @[PEArray.scala 202:32 PEArray.scala 203:15]
  wire [2:0] _GEN_331 = count == count_max ? 3'h0 : state; // @[PEArray.scala 202:32 PEArray.scala 204:15 PEArray.scala 100:22]
  wire [9:0] _GEN_865 = {{4'd0}, GRU_out_width}; // @[PEArray.scala 220:19]
  wire [9:0] _GEN_0 = count % _GEN_865; // @[PEArray.scala 220:19]
  wire [5:0] _T_36 = _GEN_0[5:0]; // @[PEArray.scala 220:19]
  wire [5:0] _T_38 = GRU_out_width - 6'h1; // @[PEArray.scala 220:55]
  wire [5:0] _GEN_334 = _T_36 == _T_38 ? _L0Index_T_2 : L0index_begin; // @[PEArray.scala 220:62 PEArray.scala 221:17 PEArray.scala 214:15]
  wire [5:0] _GEN_346 = _T_41 ? _GEN_334 : L0Index; // @[Conditional.scala 39:67 PEArray.scala 39:24]
  wire [9:0] _GEN_347 = _T_41 ? _GEN_330 : count; // @[Conditional.scala 39:67 PEArray.scala 101:22]
  wire [2:0] _GEN_348 = _T_41 ? _GEN_331 : state; // @[Conditional.scala 39:67 PEArray.scala 100:22]
  wire [5:0] _GEN_353 = _T_31 ? _GEN_334 : _GEN_346; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_354 = _T_31 ? _GEN_330 : _GEN_347; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_355 = _T_31 ? _GEN_331 : _GEN_348; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_356 = _T_22 ? _GEN_330 : _GEN_354; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_357 = _T_22 ? _GEN_329 : _GEN_353; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_458 = _T_22 ? _GEN_331 : _GEN_355; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_690 = _T_3 ? _GEN_118 : {{2'd0}, GRU_out_width}; // @[Conditional.scala 40:58 PEArray.scala 104:26]
  FP16MulAdder FP16MAC ( // @[PEArray.scala 72:23]
    .io_a(FP16MAC_io_a),
    .io_b(FP16MAC_io_b),
    .io_c(FP16MAC_io_c),
    .io_out(FP16MAC_io_out)
  );
  assign io_ToRightPE = mux3out_reg; // @[PEArray.scala 95:16]
  assign io_ToBelowPE = mux2out_reg; // @[PEArray.scala 94:16]
  assign FP16MAC_io_a = sel1 ? io_FromL1 : io_FromLeftPE; // @[PEArray.scala 50:14 PEArray.scala 50:23 PEArray.scala 51:24]
  assign FP16MAC_io_b = sel5 ? mux4out : _GEN_105; // @[PEArray.scala 77:13 PEArray.scala 78:18 PEArray.scala 81:18]
  assign FP16MAC_io_c = sel5 ? _GEN_105 : mux4out; // @[PEArray.scala 77:13 PEArray.scala 79:18 PEArray.scala 82:18]
  always @(posedge clock) begin
    if (reset) begin // @[PEArray.scala 39:24]
      L0Index <= 6'h0; // @[PEArray.scala 39:24]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h2; // @[PEArray.scala 159:15]
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h7; // @[PEArray.scala 181:15]
      end else begin
        L0Index <= _GEN_357;
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_0 <= _GEN_229;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_1 <= _GEN_230;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_2 <= _GEN_231;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_3 <= _GEN_232;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_4 <= _GEN_233;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_5 <= _GEN_234;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_6 <= _GEN_235;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_7 <= _GEN_236;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_8 <= _GEN_237;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_9 <= _GEN_238;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_10 <= _GEN_239;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_11 <= _GEN_240;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_12 <= _GEN_241;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_13 <= _GEN_242;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_14 <= _GEN_243;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_15 <= _GEN_244;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_16 <= _GEN_245;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_17 <= _GEN_246;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_18 <= _GEN_247;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_19 <= _GEN_248;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_20 <= _GEN_249;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_21 <= _GEN_250;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_22 <= _GEN_251;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_23 <= _GEN_252;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_24 <= _GEN_253;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_25 <= _GEN_254;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_26 <= _GEN_255;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_27 <= _GEN_256;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_28 <= _GEN_257;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_29 <= _GEN_258;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_30 <= _GEN_259;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_31 <= _GEN_260;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_32 <= _GEN_261;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_33 <= _GEN_262;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_34 <= _GEN_263;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_35 <= _GEN_264;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_36 <= _GEN_265;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_37 <= _GEN_266;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_38 <= _GEN_267;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_39 <= _GEN_268;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_40 <= _GEN_269;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_41 <= _GEN_270;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_42 <= _GEN_271;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_43 <= _GEN_272;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_44 <= _GEN_273;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_45 <= _GEN_274;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_46 <= _GEN_275;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_47 <= _GEN_276;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_48 <= _GEN_277;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_49 <= _GEN_278;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_50 <= _GEN_279;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_51 <= _GEN_280;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_52 <= _GEN_281;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_53 <= _GEN_282;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_54 <= _GEN_283;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_55 <= _GEN_284;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_56 <= _GEN_285;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_57 <= _GEN_286;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_58 <= _GEN_287;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_59 <= _GEN_288;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_60 <= _GEN_289;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_61 <= _GEN_290;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_62 <= _GEN_291;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_63 <= _GEN_292;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_64 <= _GEN_293;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_65 <= _GEN_294;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_66 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_67 <= _GEN_296;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_68 <= _GEN_297;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_69 <= _GEN_298;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_70 <= _GEN_299;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_71 <= _GEN_300;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_72 <= _GEN_301;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_73 <= _GEN_302;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_74 <= _GEN_303;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_75 <= _GEN_304;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_76 <= _GEN_305;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_77 <= _GEN_306;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_78 <= _GEN_307;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_79 <= _GEN_308;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_80 <= _GEN_309;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_81 <= _GEN_310;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_82 <= _GEN_311;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_83 <= _GEN_312;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_84 <= _GEN_313;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_85 <= _GEN_314;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_86 <= _GEN_315;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_87 <= _GEN_316;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_88 <= _GEN_317;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_89 <= _GEN_318;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_90 <= _GEN_319;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_91 <= _GEN_320;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_92 <= _GEN_321;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_93 <= _GEN_322;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_94 <= _GEN_323;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_95 <= _GEN_324;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_96 <= _GEN_325;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_97 <= _GEN_326;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_98 <= _GEN_327;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_99 <= _GEN_328;
          end
        end
      end
    end
    if (reset) begin // @[PEArray.scala 100:22]
      state <= 3'h0; // @[PEArray.scala 100:22]
    end else if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[7]) begin // @[PEArray.scala 116:57]
        if (_T_6) begin // @[Conditional.scala 40:58]
          state <= 3'h0; // @[PEArray.scala 120:19]
        end else begin
          state <= _GEN_113;
        end
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      if (count == 10'h33) begin // @[PEArray.scala 164:27]
        state <= 3'h0; // @[PEArray.scala 166:15]
      end
    end else if (_T_16) begin // @[Conditional.scala 39:67]
      state <= _GEN_126;
    end else begin
      state <= _GEN_458;
    end
    if (reset) begin // @[PEArray.scala 90:28]
      mux2out_reg <= 16'h0; // @[PEArray.scala 90:28]
    end else begin
      mux2out_reg <= MAC_out; // @[PEArray.scala 90:28]
    end
    if (reset) begin // @[PEArray.scala 91:28]
      mux3out_reg <= 16'h0; // @[PEArray.scala 91:28]
    end else if (sel3) begin // @[PEArray.scala 56:14]
      mux3out_reg <= MAC_out; // @[PEArray.scala 56:23]
    end else if (sel1) begin // @[PEArray.scala 50:14]
      mux3out_reg <= io_FromL1; // @[PEArray.scala 50:23]
    end else begin
      mux3out_reg <= io_FromLeftPE; // @[PEArray.scala 51:24]
    end
    if (reset) begin // @[PEArray.scala 101:22]
      count <= 10'h0; // @[PEArray.scala 101:22]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        if (count == 10'h33) begin // @[PEArray.scala 164:27]
          count <= 10'h0; // @[PEArray.scala 165:15]
        end else begin
          count <= _GEN_120;
        end
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        count <= _GEN_125;
      end else begin
        count <= _GEN_356;
      end
    end
    if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[7]) begin // @[PEArray.scala 116:57]
        count_max <= io_control_signal_count; // @[PEArray.scala 143:19]
      end
    end
    if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[7]) begin // @[PEArray.scala 116:57]
        L0index_begin <= io_control_signal_L0index; // @[PEArray.scala 144:23]
      end
    end
    GRU_out_width <= _GEN_690[5:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  L0Index = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  L0Memory_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  L0Memory_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  L0Memory_2 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  L0Memory_3 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  L0Memory_4 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  L0Memory_5 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  L0Memory_6 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  L0Memory_7 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  L0Memory_8 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  L0Memory_9 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  L0Memory_10 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  L0Memory_11 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  L0Memory_12 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  L0Memory_13 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  L0Memory_14 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  L0Memory_15 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  L0Memory_16 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  L0Memory_17 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  L0Memory_18 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  L0Memory_19 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  L0Memory_20 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  L0Memory_21 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  L0Memory_22 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  L0Memory_23 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  L0Memory_24 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  L0Memory_25 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  L0Memory_26 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  L0Memory_27 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  L0Memory_28 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  L0Memory_29 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  L0Memory_30 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  L0Memory_31 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  L0Memory_32 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  L0Memory_33 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  L0Memory_34 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  L0Memory_35 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  L0Memory_36 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  L0Memory_37 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  L0Memory_38 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  L0Memory_39 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  L0Memory_40 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  L0Memory_41 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  L0Memory_42 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  L0Memory_43 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  L0Memory_44 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  L0Memory_45 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  L0Memory_46 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  L0Memory_47 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  L0Memory_48 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  L0Memory_49 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  L0Memory_50 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  L0Memory_51 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  L0Memory_52 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  L0Memory_53 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  L0Memory_54 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  L0Memory_55 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  L0Memory_56 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  L0Memory_57 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  L0Memory_58 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  L0Memory_59 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  L0Memory_60 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  L0Memory_61 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  L0Memory_62 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  L0Memory_63 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  L0Memory_64 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  L0Memory_65 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  L0Memory_66 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  L0Memory_67 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  L0Memory_68 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  L0Memory_69 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  L0Memory_70 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  L0Memory_71 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  L0Memory_72 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  L0Memory_73 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  L0Memory_74 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  L0Memory_75 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  L0Memory_76 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  L0Memory_77 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  L0Memory_78 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  L0Memory_79 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  L0Memory_80 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  L0Memory_81 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  L0Memory_82 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  L0Memory_83 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  L0Memory_84 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  L0Memory_85 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  L0Memory_86 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  L0Memory_87 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  L0Memory_88 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  L0Memory_89 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  L0Memory_90 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  L0Memory_91 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  L0Memory_92 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  L0Memory_93 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  L0Memory_94 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  L0Memory_95 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  L0Memory_96 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  L0Memory_97 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  L0Memory_98 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  L0Memory_99 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  state = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  mux2out_reg = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  mux3out_reg = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  count = _RAND_104[9:0];
  _RAND_105 = {1{`RANDOM}};
  count_max = _RAND_105[9:0];
  _RAND_106 = {1{`RANDOM}};
  L0index_begin = _RAND_106[5:0];
  _RAND_107 = {1{`RANDOM}};
  GRU_out_width = _RAND_107[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PE_15(
  input         clock,
  input         reset,
  input  [15:0] io_FromAbovePE,
  input  [15:0] io_FromLeftPE,
  input  [15:0] io_FromL1,
  input  [11:0] io_control_signal_mask,
  output [15:0] io_ToRightPE,
  output [15:0] io_ToBelowPE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] FP16MAC_io_a; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_b; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_c; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_out; // @[PEArray.scala 72:23]
  reg [5:0] L0Index; // @[PEArray.scala 39:24]
  reg [15:0] L0Memory_0; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_1; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_2; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_3; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_4; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_5; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_6; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_7; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_8; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_9; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_10; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_11; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_12; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_13; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_14; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_15; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_16; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_17; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_18; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_19; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_20; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_21; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_22; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_23; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_24; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_25; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_26; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_27; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_28; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_29; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_30; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_31; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_32; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_33; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_34; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_35; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_36; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_37; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_38; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_39; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_40; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_41; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_42; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_43; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_44; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_45; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_46; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_47; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_48; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_49; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_50; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_51; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_52; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_53; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_54; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_55; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_56; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_57; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_58; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_59; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_60; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_61; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_62; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_63; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_64; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_65; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_66; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_67; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_68; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_69; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_70; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_71; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_72; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_73; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_74; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_75; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_76; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_77; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_78; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_79; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_80; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_81; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_82; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_83; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_84; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_85; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_86; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_87; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_88; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_89; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_90; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_91; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_92; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_93; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_94; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_95; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_96; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_97; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_98; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_99; // @[PEArray.scala 40:21]
  reg [2:0] state; // @[PEArray.scala 100:22]
  wire  _T_3 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_12 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_16 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_22 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_31 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_41 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_342 = _T_41 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 231:12 PEArray.scala 32:8]
  wire  _GEN_349 = _T_31 ? 1'h0 : _GEN_342; // @[Conditional.scala 39:67 PEArray.scala 208:12]
  wire  _GEN_459 = _T_22 | _GEN_349; // @[Conditional.scala 39:67 PEArray.scala 32:8]
  wire  _GEN_463 = _T_16 ? 1'h0 : _GEN_459; // @[Conditional.scala 39:67]
  wire  _GEN_572 = _T_12 | _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 149:12]
  wire  sel1 = _T_3 | _GEN_572; // @[Conditional.scala 40:58 PEArray.scala 108:12]
  wire [15:0] MAC_out = FP16MAC_io_out; // @[PEArray.scala 47:21 PEArray.scala 85:11]
  wire  _GEN_465 = _T_16 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 177:12]
  wire  _GEN_580 = _T_12 | _GEN_465; // @[Conditional.scala 39:67 PEArray.scala 34:8]
  wire  sel3 = _T_3 | _GEN_580; // @[Conditional.scala 40:58 PEArray.scala 110:12]
  wire [1:0] _GEN_344 = _T_41 ? 2'h2 : 2'h0; // @[Conditional.scala 39:67 PEArray.scala 233:12 PEArray.scala 35:8]
  wire [1:0] _GEN_351 = _T_31 ? 2'h2 : _GEN_344; // @[Conditional.scala 39:67 PEArray.scala 210:12]
  wire [1:0] _GEN_461 = _T_22 ? 2'h0 : _GEN_351; // @[Conditional.scala 39:67 PEArray.scala 35:8]
  wire [1:0] _GEN_466 = _T_16 ? 2'h0 : _GEN_461; // @[Conditional.scala 39:67 PEArray.scala 178:12]
  wire [1:0] _GEN_574 = _T_12 ? 2'h0 : _GEN_466; // @[Conditional.scala 39:67]
  wire [1:0] sel4 = _T_3 ? 2'h0 : _GEN_574; // @[Conditional.scala 40:58 PEArray.scala 111:12]
  wire [15:0] _GEN_3 = sel4 == 2'h2 ? io_FromL1 : 16'h0; // @[PEArray.scala 65:28 PEArray.scala 66:15 PEArray.scala 69:15]
  wire [15:0] _GEN_4 = sel4 == 2'h1 ? io_FromAbovePE : _GEN_3; // @[PEArray.scala 62:28 PEArray.scala 63:15]
  wire [15:0] mux4out = sel4 == 2'h0 ? 16'h0 : _GEN_4; // @[PEArray.scala 59:22 PEArray.scala 60:13]
  wire [15:0] _GEN_7 = 6'h1 == L0Index ? L0Memory_1 : L0Memory_0; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_8 = 6'h2 == L0Index ? L0Memory_2 : _GEN_7; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_9 = 6'h3 == L0Index ? L0Memory_3 : _GEN_8; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_10 = 6'h4 == L0Index ? L0Memory_4 : _GEN_9; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_11 = 6'h5 == L0Index ? L0Memory_5 : _GEN_10; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_12 = 6'h6 == L0Index ? L0Memory_6 : _GEN_11; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_13 = 6'h7 == L0Index ? L0Memory_7 : _GEN_12; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_14 = 6'h8 == L0Index ? L0Memory_8 : _GEN_13; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_15 = 6'h9 == L0Index ? L0Memory_9 : _GEN_14; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_16 = 6'ha == L0Index ? L0Memory_10 : _GEN_15; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_17 = 6'hb == L0Index ? L0Memory_11 : _GEN_16; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_18 = 6'hc == L0Index ? L0Memory_12 : _GEN_17; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_19 = 6'hd == L0Index ? L0Memory_13 : _GEN_18; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_20 = 6'he == L0Index ? L0Memory_14 : _GEN_19; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_21 = 6'hf == L0Index ? L0Memory_15 : _GEN_20; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_22 = 6'h10 == L0Index ? L0Memory_16 : _GEN_21; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_23 = 6'h11 == L0Index ? L0Memory_17 : _GEN_22; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_24 = 6'h12 == L0Index ? L0Memory_18 : _GEN_23; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_25 = 6'h13 == L0Index ? L0Memory_19 : _GEN_24; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_26 = 6'h14 == L0Index ? L0Memory_20 : _GEN_25; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_27 = 6'h15 == L0Index ? L0Memory_21 : _GEN_26; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_28 = 6'h16 == L0Index ? L0Memory_22 : _GEN_27; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_29 = 6'h17 == L0Index ? L0Memory_23 : _GEN_28; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_30 = 6'h18 == L0Index ? L0Memory_24 : _GEN_29; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_31 = 6'h19 == L0Index ? L0Memory_25 : _GEN_30; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_32 = 6'h1a == L0Index ? L0Memory_26 : _GEN_31; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_33 = 6'h1b == L0Index ? L0Memory_27 : _GEN_32; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_34 = 6'h1c == L0Index ? L0Memory_28 : _GEN_33; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_35 = 6'h1d == L0Index ? L0Memory_29 : _GEN_34; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_36 = 6'h1e == L0Index ? L0Memory_30 : _GEN_35; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_37 = 6'h1f == L0Index ? L0Memory_31 : _GEN_36; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_38 = 6'h20 == L0Index ? L0Memory_32 : _GEN_37; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_39 = 6'h21 == L0Index ? L0Memory_33 : _GEN_38; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_40 = 6'h22 == L0Index ? L0Memory_34 : _GEN_39; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_41 = 6'h23 == L0Index ? L0Memory_35 : _GEN_40; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_42 = 6'h24 == L0Index ? L0Memory_36 : _GEN_41; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_43 = 6'h25 == L0Index ? L0Memory_37 : _GEN_42; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_44 = 6'h26 == L0Index ? L0Memory_38 : _GEN_43; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_45 = 6'h27 == L0Index ? L0Memory_39 : _GEN_44; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_46 = 6'h28 == L0Index ? L0Memory_40 : _GEN_45; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_47 = 6'h29 == L0Index ? L0Memory_41 : _GEN_46; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_48 = 6'h2a == L0Index ? L0Memory_42 : _GEN_47; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_49 = 6'h2b == L0Index ? L0Memory_43 : _GEN_48; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_50 = 6'h2c == L0Index ? L0Memory_44 : _GEN_49; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_51 = 6'h2d == L0Index ? L0Memory_45 : _GEN_50; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_52 = 6'h2e == L0Index ? L0Memory_46 : _GEN_51; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_53 = 6'h2f == L0Index ? L0Memory_47 : _GEN_52; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_54 = 6'h30 == L0Index ? L0Memory_48 : _GEN_53; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_55 = 6'h31 == L0Index ? L0Memory_49 : _GEN_54; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_56 = 6'h32 == L0Index ? L0Memory_50 : _GEN_55; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_57 = 6'h33 == L0Index ? L0Memory_51 : _GEN_56; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_58 = 6'h34 == L0Index ? L0Memory_52 : _GEN_57; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_59 = 6'h35 == L0Index ? L0Memory_53 : _GEN_58; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_60 = 6'h36 == L0Index ? L0Memory_54 : _GEN_59; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_61 = 6'h37 == L0Index ? L0Memory_55 : _GEN_60; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_62 = 6'h38 == L0Index ? L0Memory_56 : _GEN_61; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_63 = 6'h39 == L0Index ? L0Memory_57 : _GEN_62; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_64 = 6'h3a == L0Index ? L0Memory_58 : _GEN_63; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_65 = 6'h3b == L0Index ? L0Memory_59 : _GEN_64; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_66 = 6'h3c == L0Index ? L0Memory_60 : _GEN_65; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_67 = 6'h3d == L0Index ? L0Memory_61 : _GEN_66; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_68 = 6'h3e == L0Index ? L0Memory_62 : _GEN_67; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_69 = 6'h3f == L0Index ? L0Memory_63 : _GEN_68; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [6:0] _GEN_793 = {{1'd0}, L0Index}; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_70 = 7'h40 == _GEN_793 ? L0Memory_64 : _GEN_69; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_71 = 7'h41 == _GEN_793 ? L0Memory_65 : _GEN_70; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_72 = 7'h42 == _GEN_793 ? L0Memory_66 : _GEN_71; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_73 = 7'h43 == _GEN_793 ? L0Memory_67 : _GEN_72; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_74 = 7'h44 == _GEN_793 ? L0Memory_68 : _GEN_73; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_75 = 7'h45 == _GEN_793 ? L0Memory_69 : _GEN_74; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_76 = 7'h46 == _GEN_793 ? L0Memory_70 : _GEN_75; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_77 = 7'h47 == _GEN_793 ? L0Memory_71 : _GEN_76; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_78 = 7'h48 == _GEN_793 ? L0Memory_72 : _GEN_77; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_79 = 7'h49 == _GEN_793 ? L0Memory_73 : _GEN_78; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_80 = 7'h4a == _GEN_793 ? L0Memory_74 : _GEN_79; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_81 = 7'h4b == _GEN_793 ? L0Memory_75 : _GEN_80; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_82 = 7'h4c == _GEN_793 ? L0Memory_76 : _GEN_81; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_83 = 7'h4d == _GEN_793 ? L0Memory_77 : _GEN_82; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_84 = 7'h4e == _GEN_793 ? L0Memory_78 : _GEN_83; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_85 = 7'h4f == _GEN_793 ? L0Memory_79 : _GEN_84; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_86 = 7'h50 == _GEN_793 ? L0Memory_80 : _GEN_85; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_87 = 7'h51 == _GEN_793 ? L0Memory_81 : _GEN_86; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_88 = 7'h52 == _GEN_793 ? L0Memory_82 : _GEN_87; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_89 = 7'h53 == _GEN_793 ? L0Memory_83 : _GEN_88; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_90 = 7'h54 == _GEN_793 ? L0Memory_84 : _GEN_89; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_91 = 7'h55 == _GEN_793 ? L0Memory_85 : _GEN_90; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_92 = 7'h56 == _GEN_793 ? L0Memory_86 : _GEN_91; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_93 = 7'h57 == _GEN_793 ? L0Memory_87 : _GEN_92; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_94 = 7'h58 == _GEN_793 ? L0Memory_88 : _GEN_93; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_95 = 7'h59 == _GEN_793 ? L0Memory_89 : _GEN_94; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_96 = 7'h5a == _GEN_793 ? L0Memory_90 : _GEN_95; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_97 = 7'h5b == _GEN_793 ? L0Memory_91 : _GEN_96; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_98 = 7'h5c == _GEN_793 ? L0Memory_92 : _GEN_97; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_99 = 7'h5d == _GEN_793 ? L0Memory_93 : _GEN_98; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_100 = 7'h5e == _GEN_793 ? L0Memory_94 : _GEN_99; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_101 = 7'h5f == _GEN_793 ? L0Memory_95 : _GEN_100; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_102 = 7'h60 == _GEN_793 ? L0Memory_96 : _GEN_101; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_103 = 7'h61 == _GEN_793 ? L0Memory_97 : _GEN_102; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_104 = 7'h62 == _GEN_793 ? L0Memory_98 : _GEN_103; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_105 = 7'h63 == _GEN_793 ? L0Memory_99 : _GEN_104; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire  _GEN_575 = _T_12 ? 1'h0 : _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 157:12]
  wire  sel5 = _T_3 ? 1'h0 : _GEN_575; // @[Conditional.scala 40:58 PEArray.scala 112:12]
  reg [15:0] mux2out_reg; // @[PEArray.scala 90:28]
  reg [15:0] mux3out_reg; // @[PEArray.scala 91:28]
  reg [9:0] count; // @[PEArray.scala 101:22]
  reg [5:0] GRU_out_width; // @[PEArray.scala 104:26]
  wire [7:0] _GEN_118 = io_control_signal_mask[6] ? 8'h0 : {{2'd0}, GRU_out_width}; // @[PEArray.scala 116:57 PEArray.scala 145:23 PEArray.scala 104:26]
  wire [9:0] _count_T_1 = count + 10'h1; // @[PEArray.scala 162:24]
  wire [9:0] _GEN_120 = count != 10'h33 ? _count_T_1 : count; // @[PEArray.scala 161:27 PEArray.scala 162:15 PEArray.scala 101:22]
  wire [9:0] _GEN_124 = count != 10'h188 ? _count_T_1 : count; // @[PEArray.scala 183:28 PEArray.scala 184:15 PEArray.scala 101:22]
  wire [9:0] _GEN_125 = count == 10'h188 ? 10'h0 : _GEN_124; // @[PEArray.scala 186:28 PEArray.scala 187:15]
  wire [2:0] _GEN_126 = count == 10'h188 ? 3'h0 : state; // @[PEArray.scala 186:28 PEArray.scala 188:15 PEArray.scala 100:22]
  wire [9:0] _GEN_127 = count != 10'h0 ? _count_T_1 : count; // @[PEArray.scala 192:32 PEArray.scala 193:15 PEArray.scala 101:22]
  wire  _T_24 = count == 10'h0; // @[PEArray.scala 195:18]
  wire [5:0] _GEN_128 = count == 10'h0 ? 6'h0 : L0Index; // @[PEArray.scala 195:26 PEArray.scala 196:17 PEArray.scala 39:24]
  wire [9:0] _T_27 = 10'h0 - 10'h1; // @[PEArray.scala 198:51]
  wire [15:0] _GEN_129 = 6'h0 == L0Index ? io_FromL1 : L0Memory_0; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_130 = 6'h1 == L0Index ? io_FromL1 : L0Memory_1; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_131 = 6'h2 == L0Index ? io_FromL1 : L0Memory_2; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_132 = 6'h3 == L0Index ? io_FromL1 : L0Memory_3; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_133 = 6'h4 == L0Index ? io_FromL1 : L0Memory_4; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_134 = 6'h5 == L0Index ? io_FromL1 : L0Memory_5; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_135 = 6'h6 == L0Index ? io_FromL1 : L0Memory_6; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_136 = 6'h7 == L0Index ? io_FromL1 : L0Memory_7; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_137 = 6'h8 == L0Index ? io_FromL1 : L0Memory_8; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_138 = 6'h9 == L0Index ? io_FromL1 : L0Memory_9; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_139 = 6'ha == L0Index ? io_FromL1 : L0Memory_10; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_140 = 6'hb == L0Index ? io_FromL1 : L0Memory_11; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_141 = 6'hc == L0Index ? io_FromL1 : L0Memory_12; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_142 = 6'hd == L0Index ? io_FromL1 : L0Memory_13; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_143 = 6'he == L0Index ? io_FromL1 : L0Memory_14; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_144 = 6'hf == L0Index ? io_FromL1 : L0Memory_15; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_145 = 6'h10 == L0Index ? io_FromL1 : L0Memory_16; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_146 = 6'h11 == L0Index ? io_FromL1 : L0Memory_17; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_147 = 6'h12 == L0Index ? io_FromL1 : L0Memory_18; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_148 = 6'h13 == L0Index ? io_FromL1 : L0Memory_19; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_149 = 6'h14 == L0Index ? io_FromL1 : L0Memory_20; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_150 = 6'h15 == L0Index ? io_FromL1 : L0Memory_21; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_151 = 6'h16 == L0Index ? io_FromL1 : L0Memory_22; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_152 = 6'h17 == L0Index ? io_FromL1 : L0Memory_23; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_153 = 6'h18 == L0Index ? io_FromL1 : L0Memory_24; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_154 = 6'h19 == L0Index ? io_FromL1 : L0Memory_25; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_155 = 6'h1a == L0Index ? io_FromL1 : L0Memory_26; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_156 = 6'h1b == L0Index ? io_FromL1 : L0Memory_27; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_157 = 6'h1c == L0Index ? io_FromL1 : L0Memory_28; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_158 = 6'h1d == L0Index ? io_FromL1 : L0Memory_29; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_159 = 6'h1e == L0Index ? io_FromL1 : L0Memory_30; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_160 = 6'h1f == L0Index ? io_FromL1 : L0Memory_31; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_161 = 6'h20 == L0Index ? io_FromL1 : L0Memory_32; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_162 = 6'h21 == L0Index ? io_FromL1 : L0Memory_33; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_163 = 6'h22 == L0Index ? io_FromL1 : L0Memory_34; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_164 = 6'h23 == L0Index ? io_FromL1 : L0Memory_35; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_165 = 6'h24 == L0Index ? io_FromL1 : L0Memory_36; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_166 = 6'h25 == L0Index ? io_FromL1 : L0Memory_37; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_167 = 6'h26 == L0Index ? io_FromL1 : L0Memory_38; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_168 = 6'h27 == L0Index ? io_FromL1 : L0Memory_39; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_169 = 6'h28 == L0Index ? io_FromL1 : L0Memory_40; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_170 = 6'h29 == L0Index ? io_FromL1 : L0Memory_41; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_171 = 6'h2a == L0Index ? io_FromL1 : L0Memory_42; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_172 = 6'h2b == L0Index ? io_FromL1 : L0Memory_43; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_173 = 6'h2c == L0Index ? io_FromL1 : L0Memory_44; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_174 = 6'h2d == L0Index ? io_FromL1 : L0Memory_45; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_175 = 6'h2e == L0Index ? io_FromL1 : L0Memory_46; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_176 = 6'h2f == L0Index ? io_FromL1 : L0Memory_47; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_177 = 6'h30 == L0Index ? io_FromL1 : L0Memory_48; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_178 = 6'h31 == L0Index ? io_FromL1 : L0Memory_49; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_179 = 6'h32 == L0Index ? io_FromL1 : L0Memory_50; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_180 = 6'h33 == L0Index ? io_FromL1 : L0Memory_51; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_181 = 6'h34 == L0Index ? io_FromL1 : L0Memory_52; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_182 = 6'h35 == L0Index ? io_FromL1 : L0Memory_53; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_183 = 6'h36 == L0Index ? io_FromL1 : L0Memory_54; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_184 = 6'h37 == L0Index ? io_FromL1 : L0Memory_55; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_185 = 6'h38 == L0Index ? io_FromL1 : L0Memory_56; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_186 = 6'h39 == L0Index ? io_FromL1 : L0Memory_57; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_187 = 6'h3a == L0Index ? io_FromL1 : L0Memory_58; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_188 = 6'h3b == L0Index ? io_FromL1 : L0Memory_59; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_189 = 6'h3c == L0Index ? io_FromL1 : L0Memory_60; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_190 = 6'h3d == L0Index ? io_FromL1 : L0Memory_61; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_191 = 6'h3e == L0Index ? io_FromL1 : L0Memory_62; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_192 = 6'h3f == L0Index ? io_FromL1 : L0Memory_63; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_193 = 7'h40 == _GEN_793 ? io_FromL1 : L0Memory_64; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_194 = 7'h41 == _GEN_793 ? io_FromL1 : L0Memory_65; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_195 = 7'h42 == _GEN_793 ? io_FromL1 : L0Memory_66; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_196 = 7'h43 == _GEN_793 ? io_FromL1 : L0Memory_67; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_197 = 7'h44 == _GEN_793 ? io_FromL1 : L0Memory_68; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_198 = 7'h45 == _GEN_793 ? io_FromL1 : L0Memory_69; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_199 = 7'h46 == _GEN_793 ? io_FromL1 : L0Memory_70; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_200 = 7'h47 == _GEN_793 ? io_FromL1 : L0Memory_71; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_201 = 7'h48 == _GEN_793 ? io_FromL1 : L0Memory_72; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_202 = 7'h49 == _GEN_793 ? io_FromL1 : L0Memory_73; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_203 = 7'h4a == _GEN_793 ? io_FromL1 : L0Memory_74; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_204 = 7'h4b == _GEN_793 ? io_FromL1 : L0Memory_75; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_205 = 7'h4c == _GEN_793 ? io_FromL1 : L0Memory_76; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_206 = 7'h4d == _GEN_793 ? io_FromL1 : L0Memory_77; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_207 = 7'h4e == _GEN_793 ? io_FromL1 : L0Memory_78; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_208 = 7'h4f == _GEN_793 ? io_FromL1 : L0Memory_79; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_209 = 7'h50 == _GEN_793 ? io_FromL1 : L0Memory_80; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_210 = 7'h51 == _GEN_793 ? io_FromL1 : L0Memory_81; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_211 = 7'h52 == _GEN_793 ? io_FromL1 : L0Memory_82; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_212 = 7'h53 == _GEN_793 ? io_FromL1 : L0Memory_83; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_213 = 7'h54 == _GEN_793 ? io_FromL1 : L0Memory_84; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_214 = 7'h55 == _GEN_793 ? io_FromL1 : L0Memory_85; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_215 = 7'h56 == _GEN_793 ? io_FromL1 : L0Memory_86; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_216 = 7'h57 == _GEN_793 ? io_FromL1 : L0Memory_87; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_217 = 7'h58 == _GEN_793 ? io_FromL1 : L0Memory_88; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_218 = 7'h59 == _GEN_793 ? io_FromL1 : L0Memory_89; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_219 = 7'h5a == _GEN_793 ? io_FromL1 : L0Memory_90; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_220 = 7'h5b == _GEN_793 ? io_FromL1 : L0Memory_91; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_221 = 7'h5c == _GEN_793 ? io_FromL1 : L0Memory_92; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_222 = 7'h5d == _GEN_793 ? io_FromL1 : L0Memory_93; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_223 = 7'h5e == _GEN_793 ? io_FromL1 : L0Memory_94; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_224 = 7'h5f == _GEN_793 ? io_FromL1 : L0Memory_95; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_225 = 7'h60 == _GEN_793 ? io_FromL1 : L0Memory_96; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_226 = 7'h61 == _GEN_793 ? io_FromL1 : L0Memory_97; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_227 = 7'h62 == _GEN_793 ? io_FromL1 : L0Memory_98; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_228 = 7'h63 == _GEN_793 ? io_FromL1 : L0Memory_99; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [5:0] _L0Index_T_2 = L0Index + 6'h1; // @[PEArray.scala 200:28]
  wire [15:0] _GEN_229 = count >= 10'h1 & count <= _T_27 ? _GEN_129 : L0Memory_0; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_230 = count >= 10'h1 & count <= _T_27 ? _GEN_130 : L0Memory_1; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_231 = count >= 10'h1 & count <= _T_27 ? _GEN_131 : L0Memory_2; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_232 = count >= 10'h1 & count <= _T_27 ? _GEN_132 : L0Memory_3; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_233 = count >= 10'h1 & count <= _T_27 ? _GEN_133 : L0Memory_4; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_234 = count >= 10'h1 & count <= _T_27 ? _GEN_134 : L0Memory_5; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_235 = count >= 10'h1 & count <= _T_27 ? _GEN_135 : L0Memory_6; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_236 = count >= 10'h1 & count <= _T_27 ? _GEN_136 : L0Memory_7; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_237 = count >= 10'h1 & count <= _T_27 ? _GEN_137 : L0Memory_8; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_238 = count >= 10'h1 & count <= _T_27 ? _GEN_138 : L0Memory_9; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_239 = count >= 10'h1 & count <= _T_27 ? _GEN_139 : L0Memory_10; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_240 = count >= 10'h1 & count <= _T_27 ? _GEN_140 : L0Memory_11; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_241 = count >= 10'h1 & count <= _T_27 ? _GEN_141 : L0Memory_12; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_242 = count >= 10'h1 & count <= _T_27 ? _GEN_142 : L0Memory_13; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_243 = count >= 10'h1 & count <= _T_27 ? _GEN_143 : L0Memory_14; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_244 = count >= 10'h1 & count <= _T_27 ? _GEN_144 : L0Memory_15; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_245 = count >= 10'h1 & count <= _T_27 ? _GEN_145 : L0Memory_16; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_246 = count >= 10'h1 & count <= _T_27 ? _GEN_146 : L0Memory_17; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_247 = count >= 10'h1 & count <= _T_27 ? _GEN_147 : L0Memory_18; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_248 = count >= 10'h1 & count <= _T_27 ? _GEN_148 : L0Memory_19; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_249 = count >= 10'h1 & count <= _T_27 ? _GEN_149 : L0Memory_20; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_250 = count >= 10'h1 & count <= _T_27 ? _GEN_150 : L0Memory_21; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_251 = count >= 10'h1 & count <= _T_27 ? _GEN_151 : L0Memory_22; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_252 = count >= 10'h1 & count <= _T_27 ? _GEN_152 : L0Memory_23; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_253 = count >= 10'h1 & count <= _T_27 ? _GEN_153 : L0Memory_24; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_254 = count >= 10'h1 & count <= _T_27 ? _GEN_154 : L0Memory_25; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_255 = count >= 10'h1 & count <= _T_27 ? _GEN_155 : L0Memory_26; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_256 = count >= 10'h1 & count <= _T_27 ? _GEN_156 : L0Memory_27; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_257 = count >= 10'h1 & count <= _T_27 ? _GEN_157 : L0Memory_28; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_258 = count >= 10'h1 & count <= _T_27 ? _GEN_158 : L0Memory_29; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_259 = count >= 10'h1 & count <= _T_27 ? _GEN_159 : L0Memory_30; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_260 = count >= 10'h1 & count <= _T_27 ? _GEN_160 : L0Memory_31; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_261 = count >= 10'h1 & count <= _T_27 ? _GEN_161 : L0Memory_32; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_262 = count >= 10'h1 & count <= _T_27 ? _GEN_162 : L0Memory_33; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_263 = count >= 10'h1 & count <= _T_27 ? _GEN_163 : L0Memory_34; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_264 = count >= 10'h1 & count <= _T_27 ? _GEN_164 : L0Memory_35; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_265 = count >= 10'h1 & count <= _T_27 ? _GEN_165 : L0Memory_36; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_266 = count >= 10'h1 & count <= _T_27 ? _GEN_166 : L0Memory_37; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_267 = count >= 10'h1 & count <= _T_27 ? _GEN_167 : L0Memory_38; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_268 = count >= 10'h1 & count <= _T_27 ? _GEN_168 : L0Memory_39; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_269 = count >= 10'h1 & count <= _T_27 ? _GEN_169 : L0Memory_40; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_270 = count >= 10'h1 & count <= _T_27 ? _GEN_170 : L0Memory_41; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_271 = count >= 10'h1 & count <= _T_27 ? _GEN_171 : L0Memory_42; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_272 = count >= 10'h1 & count <= _T_27 ? _GEN_172 : L0Memory_43; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_273 = count >= 10'h1 & count <= _T_27 ? _GEN_173 : L0Memory_44; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_274 = count >= 10'h1 & count <= _T_27 ? _GEN_174 : L0Memory_45; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_275 = count >= 10'h1 & count <= _T_27 ? _GEN_175 : L0Memory_46; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_276 = count >= 10'h1 & count <= _T_27 ? _GEN_176 : L0Memory_47; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_277 = count >= 10'h1 & count <= _T_27 ? _GEN_177 : L0Memory_48; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_278 = count >= 10'h1 & count <= _T_27 ? _GEN_178 : L0Memory_49; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_279 = count >= 10'h1 & count <= _T_27 ? _GEN_179 : L0Memory_50; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_280 = count >= 10'h1 & count <= _T_27 ? _GEN_180 : L0Memory_51; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_281 = count >= 10'h1 & count <= _T_27 ? _GEN_181 : L0Memory_52; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_282 = count >= 10'h1 & count <= _T_27 ? _GEN_182 : L0Memory_53; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_283 = count >= 10'h1 & count <= _T_27 ? _GEN_183 : L0Memory_54; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_284 = count >= 10'h1 & count <= _T_27 ? _GEN_184 : L0Memory_55; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_285 = count >= 10'h1 & count <= _T_27 ? _GEN_185 : L0Memory_56; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_286 = count >= 10'h1 & count <= _T_27 ? _GEN_186 : L0Memory_57; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_287 = count >= 10'h1 & count <= _T_27 ? _GEN_187 : L0Memory_58; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_288 = count >= 10'h1 & count <= _T_27 ? _GEN_188 : L0Memory_59; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_289 = count >= 10'h1 & count <= _T_27 ? _GEN_189 : L0Memory_60; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_290 = count >= 10'h1 & count <= _T_27 ? _GEN_190 : L0Memory_61; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_291 = count >= 10'h1 & count <= _T_27 ? _GEN_191 : L0Memory_62; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_292 = count >= 10'h1 & count <= _T_27 ? _GEN_192 : L0Memory_63; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_293 = count >= 10'h1 & count <= _T_27 ? _GEN_193 : L0Memory_64; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_294 = count >= 10'h1 & count <= _T_27 ? _GEN_194 : L0Memory_65; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_295 = count >= 10'h1 & count <= _T_27 ? _GEN_195 : L0Memory_66; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_296 = count >= 10'h1 & count <= _T_27 ? _GEN_196 : L0Memory_67; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_297 = count >= 10'h1 & count <= _T_27 ? _GEN_197 : L0Memory_68; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_298 = count >= 10'h1 & count <= _T_27 ? _GEN_198 : L0Memory_69; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_299 = count >= 10'h1 & count <= _T_27 ? _GEN_199 : L0Memory_70; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_300 = count >= 10'h1 & count <= _T_27 ? _GEN_200 : L0Memory_71; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_301 = count >= 10'h1 & count <= _T_27 ? _GEN_201 : L0Memory_72; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_302 = count >= 10'h1 & count <= _T_27 ? _GEN_202 : L0Memory_73; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_303 = count >= 10'h1 & count <= _T_27 ? _GEN_203 : L0Memory_74; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_304 = count >= 10'h1 & count <= _T_27 ? _GEN_204 : L0Memory_75; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_305 = count >= 10'h1 & count <= _T_27 ? _GEN_205 : L0Memory_76; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_306 = count >= 10'h1 & count <= _T_27 ? _GEN_206 : L0Memory_77; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_307 = count >= 10'h1 & count <= _T_27 ? _GEN_207 : L0Memory_78; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_308 = count >= 10'h1 & count <= _T_27 ? _GEN_208 : L0Memory_79; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_309 = count >= 10'h1 & count <= _T_27 ? _GEN_209 : L0Memory_80; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_310 = count >= 10'h1 & count <= _T_27 ? _GEN_210 : L0Memory_81; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_311 = count >= 10'h1 & count <= _T_27 ? _GEN_211 : L0Memory_82; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_312 = count >= 10'h1 & count <= _T_27 ? _GEN_212 : L0Memory_83; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_313 = count >= 10'h1 & count <= _T_27 ? _GEN_213 : L0Memory_84; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_314 = count >= 10'h1 & count <= _T_27 ? _GEN_214 : L0Memory_85; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_315 = count >= 10'h1 & count <= _T_27 ? _GEN_215 : L0Memory_86; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_316 = count >= 10'h1 & count <= _T_27 ? _GEN_216 : L0Memory_87; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_317 = count >= 10'h1 & count <= _T_27 ? _GEN_217 : L0Memory_88; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_318 = count >= 10'h1 & count <= _T_27 ? _GEN_218 : L0Memory_89; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_319 = count >= 10'h1 & count <= _T_27 ? _GEN_219 : L0Memory_90; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_320 = count >= 10'h1 & count <= _T_27 ? _GEN_220 : L0Memory_91; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_321 = count >= 10'h1 & count <= _T_27 ? _GEN_221 : L0Memory_92; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_322 = count >= 10'h1 & count <= _T_27 ? _GEN_222 : L0Memory_93; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_323 = count >= 10'h1 & count <= _T_27 ? _GEN_223 : L0Memory_94; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_324 = count >= 10'h1 & count <= _T_27 ? _GEN_224 : L0Memory_95; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_325 = count >= 10'h1 & count <= _T_27 ? _GEN_225 : L0Memory_96; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_326 = count >= 10'h1 & count <= _T_27 ? _GEN_226 : L0Memory_97; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_327 = count >= 10'h1 & count <= _T_27 ? _GEN_227 : L0Memory_98; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_328 = count >= 10'h1 & count <= _T_27 ? _GEN_228 : L0Memory_99; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [5:0] _GEN_329 = count >= 10'h1 & count <= _T_27 ? _L0Index_T_2 : _GEN_128; // @[PEArray.scala 198:59 PEArray.scala 200:17]
  wire [9:0] _GEN_330 = _T_24 ? 10'h0 : _GEN_127; // @[PEArray.scala 202:32 PEArray.scala 203:15]
  wire [2:0] _GEN_331 = _T_24 ? 3'h0 : state; // @[PEArray.scala 202:32 PEArray.scala 204:15 PEArray.scala 100:22]
  wire [9:0] _GEN_865 = {{4'd0}, GRU_out_width}; // @[PEArray.scala 220:19]
  wire [9:0] _GEN_0 = count % _GEN_865; // @[PEArray.scala 220:19]
  wire [5:0] _T_36 = _GEN_0[5:0]; // @[PEArray.scala 220:19]
  wire [5:0] _T_38 = GRU_out_width - 6'h1; // @[PEArray.scala 220:55]
  wire [5:0] _GEN_334 = _T_36 == _T_38 ? _L0Index_T_2 : 6'h0; // @[PEArray.scala 220:62 PEArray.scala 221:17 PEArray.scala 214:15]
  wire [5:0] _GEN_346 = _T_41 ? _GEN_334 : L0Index; // @[Conditional.scala 39:67 PEArray.scala 39:24]
  wire [9:0] _GEN_347 = _T_41 ? _GEN_330 : count; // @[Conditional.scala 39:67 PEArray.scala 101:22]
  wire [2:0] _GEN_348 = _T_41 ? _GEN_331 : state; // @[Conditional.scala 39:67 PEArray.scala 100:22]
  wire [5:0] _GEN_353 = _T_31 ? _GEN_334 : _GEN_346; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_354 = _T_31 ? _GEN_330 : _GEN_347; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_355 = _T_31 ? _GEN_331 : _GEN_348; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_356 = _T_22 ? _GEN_330 : _GEN_354; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_357 = _T_22 ? _GEN_329 : _GEN_353; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_458 = _T_22 ? _GEN_331 : _GEN_355; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_690 = _T_3 ? _GEN_118 : {{2'd0}, GRU_out_width}; // @[Conditional.scala 40:58 PEArray.scala 104:26]
  FP16MulAdder FP16MAC ( // @[PEArray.scala 72:23]
    .io_a(FP16MAC_io_a),
    .io_b(FP16MAC_io_b),
    .io_c(FP16MAC_io_c),
    .io_out(FP16MAC_io_out)
  );
  assign io_ToRightPE = mux3out_reg; // @[PEArray.scala 95:16]
  assign io_ToBelowPE = mux2out_reg; // @[PEArray.scala 94:16]
  assign FP16MAC_io_a = sel1 ? io_FromL1 : io_FromLeftPE; // @[PEArray.scala 50:14 PEArray.scala 50:23 PEArray.scala 51:24]
  assign FP16MAC_io_b = sel5 ? mux4out : _GEN_105; // @[PEArray.scala 77:13 PEArray.scala 78:18 PEArray.scala 81:18]
  assign FP16MAC_io_c = sel5 ? _GEN_105 : mux4out; // @[PEArray.scala 77:13 PEArray.scala 79:18 PEArray.scala 82:18]
  always @(posedge clock) begin
    if (reset) begin // @[PEArray.scala 39:24]
      L0Index <= 6'h0; // @[PEArray.scala 39:24]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h0; // @[PEArray.scala 159:15]
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h8; // @[PEArray.scala 181:15]
      end else begin
        L0Index <= _GEN_357;
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_0 <= _GEN_229;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_1 <= _GEN_230;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_2 <= _GEN_231;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_3 <= _GEN_232;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_4 <= _GEN_233;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_5 <= _GEN_234;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_6 <= _GEN_235;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_7 <= _GEN_236;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_8 <= _GEN_237;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_9 <= _GEN_238;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_10 <= _GEN_239;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_11 <= _GEN_240;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_12 <= _GEN_241;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_13 <= _GEN_242;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_14 <= _GEN_243;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_15 <= _GEN_244;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_16 <= _GEN_245;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_17 <= _GEN_246;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_18 <= _GEN_247;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_19 <= _GEN_248;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_20 <= _GEN_249;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_21 <= _GEN_250;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_22 <= _GEN_251;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_23 <= _GEN_252;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_24 <= _GEN_253;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_25 <= _GEN_254;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_26 <= _GEN_255;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_27 <= _GEN_256;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_28 <= _GEN_257;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_29 <= _GEN_258;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_30 <= _GEN_259;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_31 <= _GEN_260;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_32 <= _GEN_261;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_33 <= _GEN_262;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_34 <= _GEN_263;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_35 <= _GEN_264;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_36 <= _GEN_265;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_37 <= _GEN_266;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_38 <= _GEN_267;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_39 <= _GEN_268;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_40 <= _GEN_269;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_41 <= _GEN_270;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_42 <= _GEN_271;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_43 <= _GEN_272;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_44 <= _GEN_273;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_45 <= _GEN_274;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_46 <= _GEN_275;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_47 <= _GEN_276;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_48 <= _GEN_277;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_49 <= _GEN_278;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_50 <= _GEN_279;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_51 <= _GEN_280;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_52 <= _GEN_281;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_53 <= _GEN_282;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_54 <= _GEN_283;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_55 <= _GEN_284;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_56 <= _GEN_285;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_57 <= _GEN_286;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_58 <= _GEN_287;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_59 <= _GEN_288;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_60 <= _GEN_289;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_61 <= _GEN_290;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_62 <= _GEN_291;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_63 <= _GEN_292;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_64 <= _GEN_293;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_65 <= _GEN_294;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_66 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_67 <= _GEN_296;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_68 <= _GEN_297;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_69 <= _GEN_298;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_70 <= _GEN_299;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_71 <= _GEN_300;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_72 <= _GEN_301;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_73 <= _GEN_302;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_74 <= _GEN_303;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_75 <= _GEN_304;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_76 <= _GEN_305;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_77 <= _GEN_306;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_78 <= _GEN_307;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_79 <= _GEN_308;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_80 <= _GEN_309;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_81 <= _GEN_310;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_82 <= _GEN_311;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_83 <= _GEN_312;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_84 <= _GEN_313;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_85 <= _GEN_314;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_86 <= _GEN_315;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_87 <= _GEN_316;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_88 <= _GEN_317;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_89 <= _GEN_318;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_90 <= _GEN_319;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_91 <= _GEN_320;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_92 <= _GEN_321;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_93 <= _GEN_322;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_94 <= _GEN_323;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_95 <= _GEN_324;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_96 <= _GEN_325;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_97 <= _GEN_326;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_98 <= _GEN_327;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_99 <= _GEN_328;
          end
        end
      end
    end
    if (reset) begin // @[PEArray.scala 100:22]
      state <= 3'h0; // @[PEArray.scala 100:22]
    end else if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[6]) begin // @[PEArray.scala 116:57]
        state <= 3'h1;
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      if (count == 10'h33) begin // @[PEArray.scala 164:27]
        state <= 3'h0; // @[PEArray.scala 166:15]
      end
    end else if (_T_16) begin // @[Conditional.scala 39:67]
      state <= _GEN_126;
    end else begin
      state <= _GEN_458;
    end
    if (reset) begin // @[PEArray.scala 90:28]
      mux2out_reg <= 16'h0; // @[PEArray.scala 90:28]
    end else begin
      mux2out_reg <= MAC_out; // @[PEArray.scala 90:28]
    end
    if (reset) begin // @[PEArray.scala 91:28]
      mux3out_reg <= 16'h0; // @[PEArray.scala 91:28]
    end else if (sel3) begin // @[PEArray.scala 56:14]
      mux3out_reg <= MAC_out; // @[PEArray.scala 56:23]
    end else if (sel1) begin // @[PEArray.scala 50:14]
      mux3out_reg <= io_FromL1; // @[PEArray.scala 50:23]
    end else begin
      mux3out_reg <= io_FromLeftPE; // @[PEArray.scala 51:24]
    end
    if (reset) begin // @[PEArray.scala 101:22]
      count <= 10'h0; // @[PEArray.scala 101:22]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        if (count == 10'h33) begin // @[PEArray.scala 164:27]
          count <= 10'h0; // @[PEArray.scala 165:15]
        end else begin
          count <= _GEN_120;
        end
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        count <= _GEN_125;
      end else begin
        count <= _GEN_356;
      end
    end
    GRU_out_width <= _GEN_690[5:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  L0Index = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  L0Memory_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  L0Memory_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  L0Memory_2 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  L0Memory_3 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  L0Memory_4 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  L0Memory_5 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  L0Memory_6 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  L0Memory_7 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  L0Memory_8 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  L0Memory_9 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  L0Memory_10 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  L0Memory_11 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  L0Memory_12 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  L0Memory_13 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  L0Memory_14 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  L0Memory_15 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  L0Memory_16 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  L0Memory_17 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  L0Memory_18 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  L0Memory_19 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  L0Memory_20 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  L0Memory_21 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  L0Memory_22 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  L0Memory_23 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  L0Memory_24 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  L0Memory_25 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  L0Memory_26 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  L0Memory_27 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  L0Memory_28 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  L0Memory_29 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  L0Memory_30 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  L0Memory_31 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  L0Memory_32 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  L0Memory_33 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  L0Memory_34 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  L0Memory_35 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  L0Memory_36 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  L0Memory_37 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  L0Memory_38 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  L0Memory_39 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  L0Memory_40 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  L0Memory_41 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  L0Memory_42 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  L0Memory_43 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  L0Memory_44 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  L0Memory_45 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  L0Memory_46 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  L0Memory_47 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  L0Memory_48 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  L0Memory_49 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  L0Memory_50 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  L0Memory_51 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  L0Memory_52 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  L0Memory_53 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  L0Memory_54 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  L0Memory_55 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  L0Memory_56 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  L0Memory_57 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  L0Memory_58 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  L0Memory_59 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  L0Memory_60 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  L0Memory_61 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  L0Memory_62 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  L0Memory_63 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  L0Memory_64 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  L0Memory_65 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  L0Memory_66 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  L0Memory_67 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  L0Memory_68 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  L0Memory_69 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  L0Memory_70 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  L0Memory_71 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  L0Memory_72 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  L0Memory_73 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  L0Memory_74 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  L0Memory_75 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  L0Memory_76 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  L0Memory_77 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  L0Memory_78 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  L0Memory_79 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  L0Memory_80 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  L0Memory_81 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  L0Memory_82 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  L0Memory_83 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  L0Memory_84 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  L0Memory_85 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  L0Memory_86 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  L0Memory_87 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  L0Memory_88 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  L0Memory_89 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  L0Memory_90 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  L0Memory_91 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  L0Memory_92 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  L0Memory_93 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  L0Memory_94 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  L0Memory_95 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  L0Memory_96 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  L0Memory_97 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  L0Memory_98 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  L0Memory_99 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  state = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  mux2out_reg = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  mux3out_reg = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  count = _RAND_104[9:0];
  _RAND_105 = {1{`RANDOM}};
  GRU_out_width = _RAND_105[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PE_16(
  input         clock,
  input         reset,
  input  [15:0] io_FromAbovePE,
  input  [15:0] io_FromLeftPE,
  input  [15:0] io_FromL1,
  input  [11:0] io_control_signal_mask,
  output [15:0] io_ToRightPE,
  output [15:0] io_ToBelowPE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] FP16MAC_io_a; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_b; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_c; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_out; // @[PEArray.scala 72:23]
  reg [5:0] L0Index; // @[PEArray.scala 39:24]
  reg [15:0] L0Memory_0; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_1; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_2; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_3; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_4; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_5; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_6; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_7; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_8; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_9; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_10; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_11; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_12; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_13; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_14; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_15; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_16; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_17; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_18; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_19; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_20; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_21; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_22; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_23; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_24; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_25; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_26; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_27; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_28; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_29; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_30; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_31; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_32; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_33; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_34; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_35; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_36; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_37; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_38; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_39; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_40; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_41; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_42; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_43; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_44; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_45; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_46; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_47; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_48; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_49; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_50; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_51; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_52; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_53; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_54; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_55; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_56; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_57; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_58; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_59; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_60; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_61; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_62; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_63; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_64; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_65; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_66; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_67; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_68; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_69; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_70; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_71; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_72; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_73; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_74; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_75; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_76; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_77; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_78; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_79; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_80; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_81; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_82; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_83; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_84; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_85; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_86; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_87; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_88; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_89; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_90; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_91; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_92; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_93; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_94; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_95; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_96; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_97; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_98; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_99; // @[PEArray.scala 40:21]
  reg [2:0] state; // @[PEArray.scala 100:22]
  wire  _T_3 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_12 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_16 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_22 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_31 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_41 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_342 = _T_41 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 231:12 PEArray.scala 32:8]
  wire  _GEN_349 = _T_31 ? 1'h0 : _GEN_342; // @[Conditional.scala 39:67 PEArray.scala 208:12]
  wire  _GEN_459 = _T_22 | _GEN_349; // @[Conditional.scala 39:67 PEArray.scala 32:8]
  wire  _GEN_463 = _T_16 ? 1'h0 : _GEN_459; // @[Conditional.scala 39:67]
  wire  _GEN_572 = _T_12 | _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 149:12]
  wire  sel1 = _T_3 | _GEN_572; // @[Conditional.scala 40:58 PEArray.scala 108:12]
  wire [15:0] MAC_out = FP16MAC_io_out; // @[PEArray.scala 47:21 PEArray.scala 85:11]
  wire  _GEN_465 = _T_16 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 177:12]
  wire  _GEN_580 = _T_12 | _GEN_465; // @[Conditional.scala 39:67 PEArray.scala 34:8]
  wire  sel3 = _T_3 | _GEN_580; // @[Conditional.scala 40:58 PEArray.scala 110:12]
  wire [1:0] _GEN_344 = _T_41 ? 2'h2 : 2'h0; // @[Conditional.scala 39:67 PEArray.scala 233:12 PEArray.scala 35:8]
  wire [1:0] _GEN_351 = _T_31 ? 2'h2 : _GEN_344; // @[Conditional.scala 39:67 PEArray.scala 210:12]
  wire [1:0] _GEN_461 = _T_22 ? 2'h0 : _GEN_351; // @[Conditional.scala 39:67 PEArray.scala 35:8]
  wire [1:0] _GEN_466 = _T_16 ? 2'h0 : _GEN_461; // @[Conditional.scala 39:67 PEArray.scala 178:12]
  wire [1:0] _GEN_574 = _T_12 ? 2'h1 : _GEN_466; // @[Conditional.scala 39:67]
  wire [1:0] sel4 = _T_3 ? 2'h0 : _GEN_574; // @[Conditional.scala 40:58 PEArray.scala 111:12]
  wire [15:0] _GEN_3 = sel4 == 2'h2 ? io_FromL1 : 16'h0; // @[PEArray.scala 65:28 PEArray.scala 66:15 PEArray.scala 69:15]
  wire [15:0] _GEN_4 = sel4 == 2'h1 ? io_FromAbovePE : _GEN_3; // @[PEArray.scala 62:28 PEArray.scala 63:15]
  wire [15:0] mux4out = sel4 == 2'h0 ? 16'h0 : _GEN_4; // @[PEArray.scala 59:22 PEArray.scala 60:13]
  wire [15:0] _GEN_7 = 6'h1 == L0Index ? L0Memory_1 : L0Memory_0; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_8 = 6'h2 == L0Index ? L0Memory_2 : _GEN_7; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_9 = 6'h3 == L0Index ? L0Memory_3 : _GEN_8; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_10 = 6'h4 == L0Index ? L0Memory_4 : _GEN_9; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_11 = 6'h5 == L0Index ? L0Memory_5 : _GEN_10; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_12 = 6'h6 == L0Index ? L0Memory_6 : _GEN_11; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_13 = 6'h7 == L0Index ? L0Memory_7 : _GEN_12; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_14 = 6'h8 == L0Index ? L0Memory_8 : _GEN_13; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_15 = 6'h9 == L0Index ? L0Memory_9 : _GEN_14; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_16 = 6'ha == L0Index ? L0Memory_10 : _GEN_15; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_17 = 6'hb == L0Index ? L0Memory_11 : _GEN_16; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_18 = 6'hc == L0Index ? L0Memory_12 : _GEN_17; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_19 = 6'hd == L0Index ? L0Memory_13 : _GEN_18; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_20 = 6'he == L0Index ? L0Memory_14 : _GEN_19; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_21 = 6'hf == L0Index ? L0Memory_15 : _GEN_20; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_22 = 6'h10 == L0Index ? L0Memory_16 : _GEN_21; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_23 = 6'h11 == L0Index ? L0Memory_17 : _GEN_22; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_24 = 6'h12 == L0Index ? L0Memory_18 : _GEN_23; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_25 = 6'h13 == L0Index ? L0Memory_19 : _GEN_24; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_26 = 6'h14 == L0Index ? L0Memory_20 : _GEN_25; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_27 = 6'h15 == L0Index ? L0Memory_21 : _GEN_26; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_28 = 6'h16 == L0Index ? L0Memory_22 : _GEN_27; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_29 = 6'h17 == L0Index ? L0Memory_23 : _GEN_28; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_30 = 6'h18 == L0Index ? L0Memory_24 : _GEN_29; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_31 = 6'h19 == L0Index ? L0Memory_25 : _GEN_30; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_32 = 6'h1a == L0Index ? L0Memory_26 : _GEN_31; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_33 = 6'h1b == L0Index ? L0Memory_27 : _GEN_32; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_34 = 6'h1c == L0Index ? L0Memory_28 : _GEN_33; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_35 = 6'h1d == L0Index ? L0Memory_29 : _GEN_34; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_36 = 6'h1e == L0Index ? L0Memory_30 : _GEN_35; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_37 = 6'h1f == L0Index ? L0Memory_31 : _GEN_36; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_38 = 6'h20 == L0Index ? L0Memory_32 : _GEN_37; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_39 = 6'h21 == L0Index ? L0Memory_33 : _GEN_38; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_40 = 6'h22 == L0Index ? L0Memory_34 : _GEN_39; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_41 = 6'h23 == L0Index ? L0Memory_35 : _GEN_40; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_42 = 6'h24 == L0Index ? L0Memory_36 : _GEN_41; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_43 = 6'h25 == L0Index ? L0Memory_37 : _GEN_42; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_44 = 6'h26 == L0Index ? L0Memory_38 : _GEN_43; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_45 = 6'h27 == L0Index ? L0Memory_39 : _GEN_44; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_46 = 6'h28 == L0Index ? L0Memory_40 : _GEN_45; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_47 = 6'h29 == L0Index ? L0Memory_41 : _GEN_46; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_48 = 6'h2a == L0Index ? L0Memory_42 : _GEN_47; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_49 = 6'h2b == L0Index ? L0Memory_43 : _GEN_48; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_50 = 6'h2c == L0Index ? L0Memory_44 : _GEN_49; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_51 = 6'h2d == L0Index ? L0Memory_45 : _GEN_50; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_52 = 6'h2e == L0Index ? L0Memory_46 : _GEN_51; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_53 = 6'h2f == L0Index ? L0Memory_47 : _GEN_52; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_54 = 6'h30 == L0Index ? L0Memory_48 : _GEN_53; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_55 = 6'h31 == L0Index ? L0Memory_49 : _GEN_54; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_56 = 6'h32 == L0Index ? L0Memory_50 : _GEN_55; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_57 = 6'h33 == L0Index ? L0Memory_51 : _GEN_56; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_58 = 6'h34 == L0Index ? L0Memory_52 : _GEN_57; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_59 = 6'h35 == L0Index ? L0Memory_53 : _GEN_58; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_60 = 6'h36 == L0Index ? L0Memory_54 : _GEN_59; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_61 = 6'h37 == L0Index ? L0Memory_55 : _GEN_60; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_62 = 6'h38 == L0Index ? L0Memory_56 : _GEN_61; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_63 = 6'h39 == L0Index ? L0Memory_57 : _GEN_62; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_64 = 6'h3a == L0Index ? L0Memory_58 : _GEN_63; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_65 = 6'h3b == L0Index ? L0Memory_59 : _GEN_64; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_66 = 6'h3c == L0Index ? L0Memory_60 : _GEN_65; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_67 = 6'h3d == L0Index ? L0Memory_61 : _GEN_66; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_68 = 6'h3e == L0Index ? L0Memory_62 : _GEN_67; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_69 = 6'h3f == L0Index ? L0Memory_63 : _GEN_68; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [6:0] _GEN_793 = {{1'd0}, L0Index}; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_70 = 7'h40 == _GEN_793 ? L0Memory_64 : _GEN_69; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_71 = 7'h41 == _GEN_793 ? L0Memory_65 : _GEN_70; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_72 = 7'h42 == _GEN_793 ? L0Memory_66 : _GEN_71; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_73 = 7'h43 == _GEN_793 ? L0Memory_67 : _GEN_72; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_74 = 7'h44 == _GEN_793 ? L0Memory_68 : _GEN_73; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_75 = 7'h45 == _GEN_793 ? L0Memory_69 : _GEN_74; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_76 = 7'h46 == _GEN_793 ? L0Memory_70 : _GEN_75; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_77 = 7'h47 == _GEN_793 ? L0Memory_71 : _GEN_76; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_78 = 7'h48 == _GEN_793 ? L0Memory_72 : _GEN_77; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_79 = 7'h49 == _GEN_793 ? L0Memory_73 : _GEN_78; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_80 = 7'h4a == _GEN_793 ? L0Memory_74 : _GEN_79; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_81 = 7'h4b == _GEN_793 ? L0Memory_75 : _GEN_80; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_82 = 7'h4c == _GEN_793 ? L0Memory_76 : _GEN_81; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_83 = 7'h4d == _GEN_793 ? L0Memory_77 : _GEN_82; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_84 = 7'h4e == _GEN_793 ? L0Memory_78 : _GEN_83; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_85 = 7'h4f == _GEN_793 ? L0Memory_79 : _GEN_84; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_86 = 7'h50 == _GEN_793 ? L0Memory_80 : _GEN_85; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_87 = 7'h51 == _GEN_793 ? L0Memory_81 : _GEN_86; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_88 = 7'h52 == _GEN_793 ? L0Memory_82 : _GEN_87; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_89 = 7'h53 == _GEN_793 ? L0Memory_83 : _GEN_88; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_90 = 7'h54 == _GEN_793 ? L0Memory_84 : _GEN_89; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_91 = 7'h55 == _GEN_793 ? L0Memory_85 : _GEN_90; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_92 = 7'h56 == _GEN_793 ? L0Memory_86 : _GEN_91; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_93 = 7'h57 == _GEN_793 ? L0Memory_87 : _GEN_92; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_94 = 7'h58 == _GEN_793 ? L0Memory_88 : _GEN_93; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_95 = 7'h59 == _GEN_793 ? L0Memory_89 : _GEN_94; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_96 = 7'h5a == _GEN_793 ? L0Memory_90 : _GEN_95; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_97 = 7'h5b == _GEN_793 ? L0Memory_91 : _GEN_96; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_98 = 7'h5c == _GEN_793 ? L0Memory_92 : _GEN_97; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_99 = 7'h5d == _GEN_793 ? L0Memory_93 : _GEN_98; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_100 = 7'h5e == _GEN_793 ? L0Memory_94 : _GEN_99; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_101 = 7'h5f == _GEN_793 ? L0Memory_95 : _GEN_100; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_102 = 7'h60 == _GEN_793 ? L0Memory_96 : _GEN_101; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_103 = 7'h61 == _GEN_793 ? L0Memory_97 : _GEN_102; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_104 = 7'h62 == _GEN_793 ? L0Memory_98 : _GEN_103; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_105 = 7'h63 == _GEN_793 ? L0Memory_99 : _GEN_104; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire  _GEN_575 = _T_12 ? 1'h0 : _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 157:12]
  wire  sel5 = _T_3 ? 1'h0 : _GEN_575; // @[Conditional.scala 40:58 PEArray.scala 112:12]
  reg [15:0] mux2out_reg; // @[PEArray.scala 90:28]
  reg [15:0] mux3out_reg; // @[PEArray.scala 91:28]
  reg [9:0] count; // @[PEArray.scala 101:22]
  reg [5:0] GRU_out_width; // @[PEArray.scala 104:26]
  wire [7:0] _GEN_118 = io_control_signal_mask[6] ? 8'h0 : {{2'd0}, GRU_out_width}; // @[PEArray.scala 116:57 PEArray.scala 145:23 PEArray.scala 104:26]
  wire [9:0] _count_T_1 = count + 10'h1; // @[PEArray.scala 162:24]
  wire [9:0] _GEN_120 = count != 10'h33 ? _count_T_1 : count; // @[PEArray.scala 161:27 PEArray.scala 162:15 PEArray.scala 101:22]
  wire [9:0] _GEN_124 = count != 10'h188 ? _count_T_1 : count; // @[PEArray.scala 183:28 PEArray.scala 184:15 PEArray.scala 101:22]
  wire [9:0] _GEN_125 = count == 10'h188 ? 10'h0 : _GEN_124; // @[PEArray.scala 186:28 PEArray.scala 187:15]
  wire [2:0] _GEN_126 = count == 10'h188 ? 3'h0 : state; // @[PEArray.scala 186:28 PEArray.scala 188:15 PEArray.scala 100:22]
  wire [9:0] _GEN_127 = count != 10'h0 ? _count_T_1 : count; // @[PEArray.scala 192:32 PEArray.scala 193:15 PEArray.scala 101:22]
  wire  _T_24 = count == 10'h0; // @[PEArray.scala 195:18]
  wire [5:0] _GEN_128 = count == 10'h0 ? 6'h0 : L0Index; // @[PEArray.scala 195:26 PEArray.scala 196:17 PEArray.scala 39:24]
  wire [9:0] _T_27 = 10'h0 - 10'h1; // @[PEArray.scala 198:51]
  wire [15:0] _GEN_129 = 6'h0 == L0Index ? io_FromL1 : L0Memory_0; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_130 = 6'h1 == L0Index ? io_FromL1 : L0Memory_1; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_131 = 6'h2 == L0Index ? io_FromL1 : L0Memory_2; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_132 = 6'h3 == L0Index ? io_FromL1 : L0Memory_3; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_133 = 6'h4 == L0Index ? io_FromL1 : L0Memory_4; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_134 = 6'h5 == L0Index ? io_FromL1 : L0Memory_5; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_135 = 6'h6 == L0Index ? io_FromL1 : L0Memory_6; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_136 = 6'h7 == L0Index ? io_FromL1 : L0Memory_7; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_137 = 6'h8 == L0Index ? io_FromL1 : L0Memory_8; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_138 = 6'h9 == L0Index ? io_FromL1 : L0Memory_9; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_139 = 6'ha == L0Index ? io_FromL1 : L0Memory_10; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_140 = 6'hb == L0Index ? io_FromL1 : L0Memory_11; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_141 = 6'hc == L0Index ? io_FromL1 : L0Memory_12; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_142 = 6'hd == L0Index ? io_FromL1 : L0Memory_13; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_143 = 6'he == L0Index ? io_FromL1 : L0Memory_14; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_144 = 6'hf == L0Index ? io_FromL1 : L0Memory_15; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_145 = 6'h10 == L0Index ? io_FromL1 : L0Memory_16; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_146 = 6'h11 == L0Index ? io_FromL1 : L0Memory_17; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_147 = 6'h12 == L0Index ? io_FromL1 : L0Memory_18; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_148 = 6'h13 == L0Index ? io_FromL1 : L0Memory_19; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_149 = 6'h14 == L0Index ? io_FromL1 : L0Memory_20; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_150 = 6'h15 == L0Index ? io_FromL1 : L0Memory_21; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_151 = 6'h16 == L0Index ? io_FromL1 : L0Memory_22; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_152 = 6'h17 == L0Index ? io_FromL1 : L0Memory_23; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_153 = 6'h18 == L0Index ? io_FromL1 : L0Memory_24; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_154 = 6'h19 == L0Index ? io_FromL1 : L0Memory_25; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_155 = 6'h1a == L0Index ? io_FromL1 : L0Memory_26; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_156 = 6'h1b == L0Index ? io_FromL1 : L0Memory_27; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_157 = 6'h1c == L0Index ? io_FromL1 : L0Memory_28; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_158 = 6'h1d == L0Index ? io_FromL1 : L0Memory_29; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_159 = 6'h1e == L0Index ? io_FromL1 : L0Memory_30; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_160 = 6'h1f == L0Index ? io_FromL1 : L0Memory_31; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_161 = 6'h20 == L0Index ? io_FromL1 : L0Memory_32; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_162 = 6'h21 == L0Index ? io_FromL1 : L0Memory_33; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_163 = 6'h22 == L0Index ? io_FromL1 : L0Memory_34; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_164 = 6'h23 == L0Index ? io_FromL1 : L0Memory_35; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_165 = 6'h24 == L0Index ? io_FromL1 : L0Memory_36; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_166 = 6'h25 == L0Index ? io_FromL1 : L0Memory_37; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_167 = 6'h26 == L0Index ? io_FromL1 : L0Memory_38; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_168 = 6'h27 == L0Index ? io_FromL1 : L0Memory_39; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_169 = 6'h28 == L0Index ? io_FromL1 : L0Memory_40; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_170 = 6'h29 == L0Index ? io_FromL1 : L0Memory_41; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_171 = 6'h2a == L0Index ? io_FromL1 : L0Memory_42; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_172 = 6'h2b == L0Index ? io_FromL1 : L0Memory_43; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_173 = 6'h2c == L0Index ? io_FromL1 : L0Memory_44; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_174 = 6'h2d == L0Index ? io_FromL1 : L0Memory_45; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_175 = 6'h2e == L0Index ? io_FromL1 : L0Memory_46; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_176 = 6'h2f == L0Index ? io_FromL1 : L0Memory_47; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_177 = 6'h30 == L0Index ? io_FromL1 : L0Memory_48; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_178 = 6'h31 == L0Index ? io_FromL1 : L0Memory_49; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_179 = 6'h32 == L0Index ? io_FromL1 : L0Memory_50; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_180 = 6'h33 == L0Index ? io_FromL1 : L0Memory_51; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_181 = 6'h34 == L0Index ? io_FromL1 : L0Memory_52; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_182 = 6'h35 == L0Index ? io_FromL1 : L0Memory_53; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_183 = 6'h36 == L0Index ? io_FromL1 : L0Memory_54; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_184 = 6'h37 == L0Index ? io_FromL1 : L0Memory_55; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_185 = 6'h38 == L0Index ? io_FromL1 : L0Memory_56; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_186 = 6'h39 == L0Index ? io_FromL1 : L0Memory_57; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_187 = 6'h3a == L0Index ? io_FromL1 : L0Memory_58; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_188 = 6'h3b == L0Index ? io_FromL1 : L0Memory_59; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_189 = 6'h3c == L0Index ? io_FromL1 : L0Memory_60; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_190 = 6'h3d == L0Index ? io_FromL1 : L0Memory_61; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_191 = 6'h3e == L0Index ? io_FromL1 : L0Memory_62; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_192 = 6'h3f == L0Index ? io_FromL1 : L0Memory_63; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_193 = 7'h40 == _GEN_793 ? io_FromL1 : L0Memory_64; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_194 = 7'h41 == _GEN_793 ? io_FromL1 : L0Memory_65; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_195 = 7'h42 == _GEN_793 ? io_FromL1 : L0Memory_66; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_196 = 7'h43 == _GEN_793 ? io_FromL1 : L0Memory_67; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_197 = 7'h44 == _GEN_793 ? io_FromL1 : L0Memory_68; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_198 = 7'h45 == _GEN_793 ? io_FromL1 : L0Memory_69; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_199 = 7'h46 == _GEN_793 ? io_FromL1 : L0Memory_70; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_200 = 7'h47 == _GEN_793 ? io_FromL1 : L0Memory_71; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_201 = 7'h48 == _GEN_793 ? io_FromL1 : L0Memory_72; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_202 = 7'h49 == _GEN_793 ? io_FromL1 : L0Memory_73; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_203 = 7'h4a == _GEN_793 ? io_FromL1 : L0Memory_74; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_204 = 7'h4b == _GEN_793 ? io_FromL1 : L0Memory_75; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_205 = 7'h4c == _GEN_793 ? io_FromL1 : L0Memory_76; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_206 = 7'h4d == _GEN_793 ? io_FromL1 : L0Memory_77; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_207 = 7'h4e == _GEN_793 ? io_FromL1 : L0Memory_78; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_208 = 7'h4f == _GEN_793 ? io_FromL1 : L0Memory_79; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_209 = 7'h50 == _GEN_793 ? io_FromL1 : L0Memory_80; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_210 = 7'h51 == _GEN_793 ? io_FromL1 : L0Memory_81; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_211 = 7'h52 == _GEN_793 ? io_FromL1 : L0Memory_82; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_212 = 7'h53 == _GEN_793 ? io_FromL1 : L0Memory_83; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_213 = 7'h54 == _GEN_793 ? io_FromL1 : L0Memory_84; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_214 = 7'h55 == _GEN_793 ? io_FromL1 : L0Memory_85; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_215 = 7'h56 == _GEN_793 ? io_FromL1 : L0Memory_86; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_216 = 7'h57 == _GEN_793 ? io_FromL1 : L0Memory_87; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_217 = 7'h58 == _GEN_793 ? io_FromL1 : L0Memory_88; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_218 = 7'h59 == _GEN_793 ? io_FromL1 : L0Memory_89; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_219 = 7'h5a == _GEN_793 ? io_FromL1 : L0Memory_90; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_220 = 7'h5b == _GEN_793 ? io_FromL1 : L0Memory_91; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_221 = 7'h5c == _GEN_793 ? io_FromL1 : L0Memory_92; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_222 = 7'h5d == _GEN_793 ? io_FromL1 : L0Memory_93; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_223 = 7'h5e == _GEN_793 ? io_FromL1 : L0Memory_94; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_224 = 7'h5f == _GEN_793 ? io_FromL1 : L0Memory_95; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_225 = 7'h60 == _GEN_793 ? io_FromL1 : L0Memory_96; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_226 = 7'h61 == _GEN_793 ? io_FromL1 : L0Memory_97; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_227 = 7'h62 == _GEN_793 ? io_FromL1 : L0Memory_98; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_228 = 7'h63 == _GEN_793 ? io_FromL1 : L0Memory_99; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [5:0] _L0Index_T_2 = L0Index + 6'h1; // @[PEArray.scala 200:28]
  wire [15:0] _GEN_229 = count >= 10'h1 & count <= _T_27 ? _GEN_129 : L0Memory_0; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_230 = count >= 10'h1 & count <= _T_27 ? _GEN_130 : L0Memory_1; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_231 = count >= 10'h1 & count <= _T_27 ? _GEN_131 : L0Memory_2; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_232 = count >= 10'h1 & count <= _T_27 ? _GEN_132 : L0Memory_3; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_233 = count >= 10'h1 & count <= _T_27 ? _GEN_133 : L0Memory_4; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_234 = count >= 10'h1 & count <= _T_27 ? _GEN_134 : L0Memory_5; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_235 = count >= 10'h1 & count <= _T_27 ? _GEN_135 : L0Memory_6; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_236 = count >= 10'h1 & count <= _T_27 ? _GEN_136 : L0Memory_7; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_237 = count >= 10'h1 & count <= _T_27 ? _GEN_137 : L0Memory_8; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_238 = count >= 10'h1 & count <= _T_27 ? _GEN_138 : L0Memory_9; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_239 = count >= 10'h1 & count <= _T_27 ? _GEN_139 : L0Memory_10; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_240 = count >= 10'h1 & count <= _T_27 ? _GEN_140 : L0Memory_11; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_241 = count >= 10'h1 & count <= _T_27 ? _GEN_141 : L0Memory_12; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_242 = count >= 10'h1 & count <= _T_27 ? _GEN_142 : L0Memory_13; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_243 = count >= 10'h1 & count <= _T_27 ? _GEN_143 : L0Memory_14; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_244 = count >= 10'h1 & count <= _T_27 ? _GEN_144 : L0Memory_15; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_245 = count >= 10'h1 & count <= _T_27 ? _GEN_145 : L0Memory_16; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_246 = count >= 10'h1 & count <= _T_27 ? _GEN_146 : L0Memory_17; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_247 = count >= 10'h1 & count <= _T_27 ? _GEN_147 : L0Memory_18; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_248 = count >= 10'h1 & count <= _T_27 ? _GEN_148 : L0Memory_19; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_249 = count >= 10'h1 & count <= _T_27 ? _GEN_149 : L0Memory_20; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_250 = count >= 10'h1 & count <= _T_27 ? _GEN_150 : L0Memory_21; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_251 = count >= 10'h1 & count <= _T_27 ? _GEN_151 : L0Memory_22; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_252 = count >= 10'h1 & count <= _T_27 ? _GEN_152 : L0Memory_23; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_253 = count >= 10'h1 & count <= _T_27 ? _GEN_153 : L0Memory_24; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_254 = count >= 10'h1 & count <= _T_27 ? _GEN_154 : L0Memory_25; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_255 = count >= 10'h1 & count <= _T_27 ? _GEN_155 : L0Memory_26; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_256 = count >= 10'h1 & count <= _T_27 ? _GEN_156 : L0Memory_27; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_257 = count >= 10'h1 & count <= _T_27 ? _GEN_157 : L0Memory_28; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_258 = count >= 10'h1 & count <= _T_27 ? _GEN_158 : L0Memory_29; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_259 = count >= 10'h1 & count <= _T_27 ? _GEN_159 : L0Memory_30; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_260 = count >= 10'h1 & count <= _T_27 ? _GEN_160 : L0Memory_31; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_261 = count >= 10'h1 & count <= _T_27 ? _GEN_161 : L0Memory_32; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_262 = count >= 10'h1 & count <= _T_27 ? _GEN_162 : L0Memory_33; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_263 = count >= 10'h1 & count <= _T_27 ? _GEN_163 : L0Memory_34; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_264 = count >= 10'h1 & count <= _T_27 ? _GEN_164 : L0Memory_35; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_265 = count >= 10'h1 & count <= _T_27 ? _GEN_165 : L0Memory_36; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_266 = count >= 10'h1 & count <= _T_27 ? _GEN_166 : L0Memory_37; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_267 = count >= 10'h1 & count <= _T_27 ? _GEN_167 : L0Memory_38; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_268 = count >= 10'h1 & count <= _T_27 ? _GEN_168 : L0Memory_39; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_269 = count >= 10'h1 & count <= _T_27 ? _GEN_169 : L0Memory_40; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_270 = count >= 10'h1 & count <= _T_27 ? _GEN_170 : L0Memory_41; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_271 = count >= 10'h1 & count <= _T_27 ? _GEN_171 : L0Memory_42; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_272 = count >= 10'h1 & count <= _T_27 ? _GEN_172 : L0Memory_43; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_273 = count >= 10'h1 & count <= _T_27 ? _GEN_173 : L0Memory_44; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_274 = count >= 10'h1 & count <= _T_27 ? _GEN_174 : L0Memory_45; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_275 = count >= 10'h1 & count <= _T_27 ? _GEN_175 : L0Memory_46; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_276 = count >= 10'h1 & count <= _T_27 ? _GEN_176 : L0Memory_47; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_277 = count >= 10'h1 & count <= _T_27 ? _GEN_177 : L0Memory_48; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_278 = count >= 10'h1 & count <= _T_27 ? _GEN_178 : L0Memory_49; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_279 = count >= 10'h1 & count <= _T_27 ? _GEN_179 : L0Memory_50; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_280 = count >= 10'h1 & count <= _T_27 ? _GEN_180 : L0Memory_51; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_281 = count >= 10'h1 & count <= _T_27 ? _GEN_181 : L0Memory_52; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_282 = count >= 10'h1 & count <= _T_27 ? _GEN_182 : L0Memory_53; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_283 = count >= 10'h1 & count <= _T_27 ? _GEN_183 : L0Memory_54; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_284 = count >= 10'h1 & count <= _T_27 ? _GEN_184 : L0Memory_55; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_285 = count >= 10'h1 & count <= _T_27 ? _GEN_185 : L0Memory_56; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_286 = count >= 10'h1 & count <= _T_27 ? _GEN_186 : L0Memory_57; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_287 = count >= 10'h1 & count <= _T_27 ? _GEN_187 : L0Memory_58; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_288 = count >= 10'h1 & count <= _T_27 ? _GEN_188 : L0Memory_59; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_289 = count >= 10'h1 & count <= _T_27 ? _GEN_189 : L0Memory_60; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_290 = count >= 10'h1 & count <= _T_27 ? _GEN_190 : L0Memory_61; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_291 = count >= 10'h1 & count <= _T_27 ? _GEN_191 : L0Memory_62; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_292 = count >= 10'h1 & count <= _T_27 ? _GEN_192 : L0Memory_63; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_293 = count >= 10'h1 & count <= _T_27 ? _GEN_193 : L0Memory_64; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_294 = count >= 10'h1 & count <= _T_27 ? _GEN_194 : L0Memory_65; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_295 = count >= 10'h1 & count <= _T_27 ? _GEN_195 : L0Memory_66; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_296 = count >= 10'h1 & count <= _T_27 ? _GEN_196 : L0Memory_67; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_297 = count >= 10'h1 & count <= _T_27 ? _GEN_197 : L0Memory_68; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_298 = count >= 10'h1 & count <= _T_27 ? _GEN_198 : L0Memory_69; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_299 = count >= 10'h1 & count <= _T_27 ? _GEN_199 : L0Memory_70; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_300 = count >= 10'h1 & count <= _T_27 ? _GEN_200 : L0Memory_71; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_301 = count >= 10'h1 & count <= _T_27 ? _GEN_201 : L0Memory_72; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_302 = count >= 10'h1 & count <= _T_27 ? _GEN_202 : L0Memory_73; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_303 = count >= 10'h1 & count <= _T_27 ? _GEN_203 : L0Memory_74; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_304 = count >= 10'h1 & count <= _T_27 ? _GEN_204 : L0Memory_75; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_305 = count >= 10'h1 & count <= _T_27 ? _GEN_205 : L0Memory_76; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_306 = count >= 10'h1 & count <= _T_27 ? _GEN_206 : L0Memory_77; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_307 = count >= 10'h1 & count <= _T_27 ? _GEN_207 : L0Memory_78; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_308 = count >= 10'h1 & count <= _T_27 ? _GEN_208 : L0Memory_79; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_309 = count >= 10'h1 & count <= _T_27 ? _GEN_209 : L0Memory_80; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_310 = count >= 10'h1 & count <= _T_27 ? _GEN_210 : L0Memory_81; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_311 = count >= 10'h1 & count <= _T_27 ? _GEN_211 : L0Memory_82; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_312 = count >= 10'h1 & count <= _T_27 ? _GEN_212 : L0Memory_83; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_313 = count >= 10'h1 & count <= _T_27 ? _GEN_213 : L0Memory_84; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_314 = count >= 10'h1 & count <= _T_27 ? _GEN_214 : L0Memory_85; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_315 = count >= 10'h1 & count <= _T_27 ? _GEN_215 : L0Memory_86; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_316 = count >= 10'h1 & count <= _T_27 ? _GEN_216 : L0Memory_87; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_317 = count >= 10'h1 & count <= _T_27 ? _GEN_217 : L0Memory_88; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_318 = count >= 10'h1 & count <= _T_27 ? _GEN_218 : L0Memory_89; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_319 = count >= 10'h1 & count <= _T_27 ? _GEN_219 : L0Memory_90; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_320 = count >= 10'h1 & count <= _T_27 ? _GEN_220 : L0Memory_91; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_321 = count >= 10'h1 & count <= _T_27 ? _GEN_221 : L0Memory_92; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_322 = count >= 10'h1 & count <= _T_27 ? _GEN_222 : L0Memory_93; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_323 = count >= 10'h1 & count <= _T_27 ? _GEN_223 : L0Memory_94; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_324 = count >= 10'h1 & count <= _T_27 ? _GEN_224 : L0Memory_95; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_325 = count >= 10'h1 & count <= _T_27 ? _GEN_225 : L0Memory_96; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_326 = count >= 10'h1 & count <= _T_27 ? _GEN_226 : L0Memory_97; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_327 = count >= 10'h1 & count <= _T_27 ? _GEN_227 : L0Memory_98; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_328 = count >= 10'h1 & count <= _T_27 ? _GEN_228 : L0Memory_99; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [5:0] _GEN_329 = count >= 10'h1 & count <= _T_27 ? _L0Index_T_2 : _GEN_128; // @[PEArray.scala 198:59 PEArray.scala 200:17]
  wire [9:0] _GEN_330 = _T_24 ? 10'h0 : _GEN_127; // @[PEArray.scala 202:32 PEArray.scala 203:15]
  wire [2:0] _GEN_331 = _T_24 ? 3'h0 : state; // @[PEArray.scala 202:32 PEArray.scala 204:15 PEArray.scala 100:22]
  wire [9:0] _GEN_865 = {{4'd0}, GRU_out_width}; // @[PEArray.scala 220:19]
  wire [9:0] _GEN_0 = count % _GEN_865; // @[PEArray.scala 220:19]
  wire [5:0] _T_36 = _GEN_0[5:0]; // @[PEArray.scala 220:19]
  wire [5:0] _T_38 = GRU_out_width - 6'h1; // @[PEArray.scala 220:55]
  wire [5:0] _GEN_334 = _T_36 == _T_38 ? _L0Index_T_2 : 6'h0; // @[PEArray.scala 220:62 PEArray.scala 221:17 PEArray.scala 214:15]
  wire [5:0] _GEN_346 = _T_41 ? _GEN_334 : L0Index; // @[Conditional.scala 39:67 PEArray.scala 39:24]
  wire [9:0] _GEN_347 = _T_41 ? _GEN_330 : count; // @[Conditional.scala 39:67 PEArray.scala 101:22]
  wire [2:0] _GEN_348 = _T_41 ? _GEN_331 : state; // @[Conditional.scala 39:67 PEArray.scala 100:22]
  wire [5:0] _GEN_353 = _T_31 ? _GEN_334 : _GEN_346; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_354 = _T_31 ? _GEN_330 : _GEN_347; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_355 = _T_31 ? _GEN_331 : _GEN_348; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_356 = _T_22 ? _GEN_330 : _GEN_354; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_357 = _T_22 ? _GEN_329 : _GEN_353; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_458 = _T_22 ? _GEN_331 : _GEN_355; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_690 = _T_3 ? _GEN_118 : {{2'd0}, GRU_out_width}; // @[Conditional.scala 40:58 PEArray.scala 104:26]
  FP16MulAdder FP16MAC ( // @[PEArray.scala 72:23]
    .io_a(FP16MAC_io_a),
    .io_b(FP16MAC_io_b),
    .io_c(FP16MAC_io_c),
    .io_out(FP16MAC_io_out)
  );
  assign io_ToRightPE = mux3out_reg; // @[PEArray.scala 95:16]
  assign io_ToBelowPE = mux2out_reg; // @[PEArray.scala 94:16]
  assign FP16MAC_io_a = sel1 ? io_FromL1 : io_FromLeftPE; // @[PEArray.scala 50:14 PEArray.scala 50:23 PEArray.scala 51:24]
  assign FP16MAC_io_b = sel5 ? mux4out : _GEN_105; // @[PEArray.scala 77:13 PEArray.scala 78:18 PEArray.scala 81:18]
  assign FP16MAC_io_c = sel5 ? _GEN_105 : mux4out; // @[PEArray.scala 77:13 PEArray.scala 79:18 PEArray.scala 82:18]
  always @(posedge clock) begin
    if (reset) begin // @[PEArray.scala 39:24]
      L0Index <= 6'h0; // @[PEArray.scala 39:24]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h1; // @[PEArray.scala 159:15]
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h8; // @[PEArray.scala 181:15]
      end else begin
        L0Index <= _GEN_357;
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_0 <= _GEN_229;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_1 <= _GEN_230;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_2 <= _GEN_231;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_3 <= _GEN_232;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_4 <= _GEN_233;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_5 <= _GEN_234;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_6 <= _GEN_235;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_7 <= _GEN_236;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_8 <= _GEN_237;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_9 <= _GEN_238;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_10 <= _GEN_239;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_11 <= _GEN_240;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_12 <= _GEN_241;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_13 <= _GEN_242;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_14 <= _GEN_243;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_15 <= _GEN_244;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_16 <= _GEN_245;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_17 <= _GEN_246;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_18 <= _GEN_247;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_19 <= _GEN_248;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_20 <= _GEN_249;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_21 <= _GEN_250;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_22 <= _GEN_251;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_23 <= _GEN_252;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_24 <= _GEN_253;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_25 <= _GEN_254;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_26 <= _GEN_255;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_27 <= _GEN_256;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_28 <= _GEN_257;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_29 <= _GEN_258;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_30 <= _GEN_259;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_31 <= _GEN_260;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_32 <= _GEN_261;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_33 <= _GEN_262;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_34 <= _GEN_263;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_35 <= _GEN_264;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_36 <= _GEN_265;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_37 <= _GEN_266;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_38 <= _GEN_267;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_39 <= _GEN_268;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_40 <= _GEN_269;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_41 <= _GEN_270;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_42 <= _GEN_271;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_43 <= _GEN_272;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_44 <= _GEN_273;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_45 <= _GEN_274;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_46 <= _GEN_275;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_47 <= _GEN_276;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_48 <= _GEN_277;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_49 <= _GEN_278;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_50 <= _GEN_279;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_51 <= _GEN_280;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_52 <= _GEN_281;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_53 <= _GEN_282;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_54 <= _GEN_283;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_55 <= _GEN_284;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_56 <= _GEN_285;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_57 <= _GEN_286;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_58 <= _GEN_287;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_59 <= _GEN_288;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_60 <= _GEN_289;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_61 <= _GEN_290;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_62 <= _GEN_291;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_63 <= _GEN_292;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_64 <= _GEN_293;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_65 <= _GEN_294;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_66 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_67 <= _GEN_296;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_68 <= _GEN_297;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_69 <= _GEN_298;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_70 <= _GEN_299;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_71 <= _GEN_300;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_72 <= _GEN_301;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_73 <= _GEN_302;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_74 <= _GEN_303;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_75 <= _GEN_304;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_76 <= _GEN_305;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_77 <= _GEN_306;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_78 <= _GEN_307;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_79 <= _GEN_308;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_80 <= _GEN_309;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_81 <= _GEN_310;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_82 <= _GEN_311;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_83 <= _GEN_312;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_84 <= _GEN_313;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_85 <= _GEN_314;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_86 <= _GEN_315;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_87 <= _GEN_316;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_88 <= _GEN_317;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_89 <= _GEN_318;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_90 <= _GEN_319;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_91 <= _GEN_320;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_92 <= _GEN_321;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_93 <= _GEN_322;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_94 <= _GEN_323;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_95 <= _GEN_324;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_96 <= _GEN_325;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_97 <= _GEN_326;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_98 <= _GEN_327;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_99 <= _GEN_328;
          end
        end
      end
    end
    if (reset) begin // @[PEArray.scala 100:22]
      state <= 3'h0; // @[PEArray.scala 100:22]
    end else if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[6]) begin // @[PEArray.scala 116:57]
        state <= 3'h1;
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      if (count == 10'h33) begin // @[PEArray.scala 164:27]
        state <= 3'h0; // @[PEArray.scala 166:15]
      end
    end else if (_T_16) begin // @[Conditional.scala 39:67]
      state <= _GEN_126;
    end else begin
      state <= _GEN_458;
    end
    if (reset) begin // @[PEArray.scala 90:28]
      mux2out_reg <= 16'h0; // @[PEArray.scala 90:28]
    end else begin
      mux2out_reg <= MAC_out; // @[PEArray.scala 90:28]
    end
    if (reset) begin // @[PEArray.scala 91:28]
      mux3out_reg <= 16'h0; // @[PEArray.scala 91:28]
    end else if (sel3) begin // @[PEArray.scala 56:14]
      mux3out_reg <= MAC_out; // @[PEArray.scala 56:23]
    end else if (sel1) begin // @[PEArray.scala 50:14]
      mux3out_reg <= io_FromL1; // @[PEArray.scala 50:23]
    end else begin
      mux3out_reg <= io_FromLeftPE; // @[PEArray.scala 51:24]
    end
    if (reset) begin // @[PEArray.scala 101:22]
      count <= 10'h0; // @[PEArray.scala 101:22]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        if (count == 10'h33) begin // @[PEArray.scala 164:27]
          count <= 10'h0; // @[PEArray.scala 165:15]
        end else begin
          count <= _GEN_120;
        end
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        count <= _GEN_125;
      end else begin
        count <= _GEN_356;
      end
    end
    GRU_out_width <= _GEN_690[5:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  L0Index = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  L0Memory_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  L0Memory_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  L0Memory_2 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  L0Memory_3 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  L0Memory_4 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  L0Memory_5 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  L0Memory_6 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  L0Memory_7 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  L0Memory_8 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  L0Memory_9 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  L0Memory_10 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  L0Memory_11 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  L0Memory_12 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  L0Memory_13 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  L0Memory_14 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  L0Memory_15 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  L0Memory_16 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  L0Memory_17 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  L0Memory_18 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  L0Memory_19 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  L0Memory_20 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  L0Memory_21 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  L0Memory_22 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  L0Memory_23 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  L0Memory_24 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  L0Memory_25 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  L0Memory_26 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  L0Memory_27 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  L0Memory_28 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  L0Memory_29 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  L0Memory_30 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  L0Memory_31 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  L0Memory_32 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  L0Memory_33 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  L0Memory_34 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  L0Memory_35 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  L0Memory_36 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  L0Memory_37 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  L0Memory_38 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  L0Memory_39 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  L0Memory_40 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  L0Memory_41 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  L0Memory_42 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  L0Memory_43 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  L0Memory_44 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  L0Memory_45 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  L0Memory_46 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  L0Memory_47 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  L0Memory_48 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  L0Memory_49 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  L0Memory_50 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  L0Memory_51 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  L0Memory_52 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  L0Memory_53 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  L0Memory_54 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  L0Memory_55 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  L0Memory_56 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  L0Memory_57 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  L0Memory_58 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  L0Memory_59 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  L0Memory_60 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  L0Memory_61 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  L0Memory_62 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  L0Memory_63 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  L0Memory_64 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  L0Memory_65 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  L0Memory_66 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  L0Memory_67 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  L0Memory_68 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  L0Memory_69 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  L0Memory_70 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  L0Memory_71 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  L0Memory_72 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  L0Memory_73 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  L0Memory_74 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  L0Memory_75 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  L0Memory_76 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  L0Memory_77 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  L0Memory_78 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  L0Memory_79 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  L0Memory_80 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  L0Memory_81 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  L0Memory_82 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  L0Memory_83 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  L0Memory_84 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  L0Memory_85 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  L0Memory_86 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  L0Memory_87 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  L0Memory_88 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  L0Memory_89 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  L0Memory_90 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  L0Memory_91 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  L0Memory_92 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  L0Memory_93 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  L0Memory_94 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  L0Memory_95 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  L0Memory_96 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  L0Memory_97 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  L0Memory_98 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  L0Memory_99 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  state = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  mux2out_reg = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  mux3out_reg = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  count = _RAND_104[9:0];
  _RAND_105 = {1{`RANDOM}};
  GRU_out_width = _RAND_105[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PE_17(
  input         clock,
  input         reset,
  input  [15:0] io_FromAbovePE,
  input  [15:0] io_FromLeftPE,
  input  [15:0] io_FromL1,
  input  [2:0]  io_control_signal_control,
  input  [9:0]  io_control_signal_count,
  input  [5:0]  io_control_signal_L0index,
  input  [11:0] io_control_signal_mask,
  input  [7:0]  io_control_signal_gru_out_width,
  output [15:0] io_ToRightPE,
  output [15:0] io_ToBelowPE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] FP16MAC_io_a; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_b; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_c; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_out; // @[PEArray.scala 72:23]
  reg [5:0] L0Index; // @[PEArray.scala 39:24]
  reg [15:0] L0Memory_0; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_1; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_2; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_3; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_4; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_5; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_6; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_7; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_8; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_9; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_10; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_11; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_12; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_13; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_14; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_15; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_16; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_17; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_18; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_19; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_20; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_21; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_22; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_23; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_24; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_25; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_26; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_27; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_28; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_29; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_30; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_31; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_32; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_33; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_34; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_35; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_36; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_37; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_38; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_39; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_40; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_41; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_42; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_43; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_44; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_45; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_46; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_47; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_48; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_49; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_50; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_51; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_52; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_53; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_54; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_55; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_56; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_57; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_58; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_59; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_60; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_61; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_62; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_63; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_64; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_65; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_66; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_67; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_68; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_69; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_70; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_71; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_72; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_73; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_74; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_75; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_76; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_77; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_78; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_79; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_80; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_81; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_82; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_83; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_84; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_85; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_86; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_87; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_88; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_89; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_90; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_91; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_92; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_93; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_94; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_95; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_96; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_97; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_98; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_99; // @[PEArray.scala 40:21]
  reg [2:0] state; // @[PEArray.scala 100:22]
  wire  _T_3 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_12 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_16 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_22 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_31 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_41 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_342 = _T_41 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 231:12 PEArray.scala 32:8]
  wire  _GEN_349 = _T_31 ? 1'h0 : _GEN_342; // @[Conditional.scala 39:67 PEArray.scala 208:12]
  wire  _GEN_459 = _T_22 | _GEN_349; // @[Conditional.scala 39:67 PEArray.scala 32:8]
  wire  _GEN_463 = _T_16 ? 1'h0 : _GEN_459; // @[Conditional.scala 39:67]
  wire  _GEN_572 = _T_12 | _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 149:12]
  wire  sel1 = _T_3 | _GEN_572; // @[Conditional.scala 40:58 PEArray.scala 108:12]
  wire [15:0] MAC_out = FP16MAC_io_out; // @[PEArray.scala 47:21 PEArray.scala 85:11]
  wire  _GEN_465 = _T_16 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 177:12]
  wire  _GEN_580 = _T_12 | _GEN_465; // @[Conditional.scala 39:67 PEArray.scala 34:8]
  wire  sel3 = _T_3 | _GEN_580; // @[Conditional.scala 40:58 PEArray.scala 110:12]
  wire [1:0] _GEN_344 = _T_41 ? 2'h2 : 2'h0; // @[Conditional.scala 39:67 PEArray.scala 233:12 PEArray.scala 35:8]
  wire [1:0] _GEN_351 = _T_31 ? 2'h2 : _GEN_344; // @[Conditional.scala 39:67 PEArray.scala 210:12]
  wire [1:0] _GEN_461 = _T_22 ? 2'h0 : _GEN_351; // @[Conditional.scala 39:67 PEArray.scala 35:8]
  wire [1:0] _GEN_466 = _T_16 ? 2'h0 : _GEN_461; // @[Conditional.scala 39:67 PEArray.scala 178:12]
  wire [1:0] _GEN_574 = _T_12 ? 2'h1 : _GEN_466; // @[Conditional.scala 39:67]
  wire [1:0] sel4 = _T_3 ? 2'h0 : _GEN_574; // @[Conditional.scala 40:58 PEArray.scala 111:12]
  wire [15:0] _GEN_3 = sel4 == 2'h2 ? io_FromL1 : 16'h0; // @[PEArray.scala 65:28 PEArray.scala 66:15 PEArray.scala 69:15]
  wire [15:0] _GEN_4 = sel4 == 2'h1 ? io_FromAbovePE : _GEN_3; // @[PEArray.scala 62:28 PEArray.scala 63:15]
  wire [15:0] mux4out = sel4 == 2'h0 ? 16'h0 : _GEN_4; // @[PEArray.scala 59:22 PEArray.scala 60:13]
  wire [15:0] _GEN_7 = 6'h1 == L0Index ? L0Memory_1 : L0Memory_0; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_8 = 6'h2 == L0Index ? L0Memory_2 : _GEN_7; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_9 = 6'h3 == L0Index ? L0Memory_3 : _GEN_8; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_10 = 6'h4 == L0Index ? L0Memory_4 : _GEN_9; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_11 = 6'h5 == L0Index ? L0Memory_5 : _GEN_10; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_12 = 6'h6 == L0Index ? L0Memory_6 : _GEN_11; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_13 = 6'h7 == L0Index ? L0Memory_7 : _GEN_12; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_14 = 6'h8 == L0Index ? L0Memory_8 : _GEN_13; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_15 = 6'h9 == L0Index ? L0Memory_9 : _GEN_14; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_16 = 6'ha == L0Index ? L0Memory_10 : _GEN_15; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_17 = 6'hb == L0Index ? L0Memory_11 : _GEN_16; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_18 = 6'hc == L0Index ? L0Memory_12 : _GEN_17; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_19 = 6'hd == L0Index ? L0Memory_13 : _GEN_18; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_20 = 6'he == L0Index ? L0Memory_14 : _GEN_19; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_21 = 6'hf == L0Index ? L0Memory_15 : _GEN_20; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_22 = 6'h10 == L0Index ? L0Memory_16 : _GEN_21; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_23 = 6'h11 == L0Index ? L0Memory_17 : _GEN_22; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_24 = 6'h12 == L0Index ? L0Memory_18 : _GEN_23; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_25 = 6'h13 == L0Index ? L0Memory_19 : _GEN_24; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_26 = 6'h14 == L0Index ? L0Memory_20 : _GEN_25; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_27 = 6'h15 == L0Index ? L0Memory_21 : _GEN_26; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_28 = 6'h16 == L0Index ? L0Memory_22 : _GEN_27; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_29 = 6'h17 == L0Index ? L0Memory_23 : _GEN_28; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_30 = 6'h18 == L0Index ? L0Memory_24 : _GEN_29; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_31 = 6'h19 == L0Index ? L0Memory_25 : _GEN_30; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_32 = 6'h1a == L0Index ? L0Memory_26 : _GEN_31; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_33 = 6'h1b == L0Index ? L0Memory_27 : _GEN_32; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_34 = 6'h1c == L0Index ? L0Memory_28 : _GEN_33; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_35 = 6'h1d == L0Index ? L0Memory_29 : _GEN_34; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_36 = 6'h1e == L0Index ? L0Memory_30 : _GEN_35; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_37 = 6'h1f == L0Index ? L0Memory_31 : _GEN_36; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_38 = 6'h20 == L0Index ? L0Memory_32 : _GEN_37; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_39 = 6'h21 == L0Index ? L0Memory_33 : _GEN_38; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_40 = 6'h22 == L0Index ? L0Memory_34 : _GEN_39; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_41 = 6'h23 == L0Index ? L0Memory_35 : _GEN_40; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_42 = 6'h24 == L0Index ? L0Memory_36 : _GEN_41; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_43 = 6'h25 == L0Index ? L0Memory_37 : _GEN_42; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_44 = 6'h26 == L0Index ? L0Memory_38 : _GEN_43; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_45 = 6'h27 == L0Index ? L0Memory_39 : _GEN_44; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_46 = 6'h28 == L0Index ? L0Memory_40 : _GEN_45; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_47 = 6'h29 == L0Index ? L0Memory_41 : _GEN_46; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_48 = 6'h2a == L0Index ? L0Memory_42 : _GEN_47; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_49 = 6'h2b == L0Index ? L0Memory_43 : _GEN_48; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_50 = 6'h2c == L0Index ? L0Memory_44 : _GEN_49; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_51 = 6'h2d == L0Index ? L0Memory_45 : _GEN_50; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_52 = 6'h2e == L0Index ? L0Memory_46 : _GEN_51; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_53 = 6'h2f == L0Index ? L0Memory_47 : _GEN_52; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_54 = 6'h30 == L0Index ? L0Memory_48 : _GEN_53; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_55 = 6'h31 == L0Index ? L0Memory_49 : _GEN_54; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_56 = 6'h32 == L0Index ? L0Memory_50 : _GEN_55; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_57 = 6'h33 == L0Index ? L0Memory_51 : _GEN_56; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_58 = 6'h34 == L0Index ? L0Memory_52 : _GEN_57; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_59 = 6'h35 == L0Index ? L0Memory_53 : _GEN_58; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_60 = 6'h36 == L0Index ? L0Memory_54 : _GEN_59; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_61 = 6'h37 == L0Index ? L0Memory_55 : _GEN_60; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_62 = 6'h38 == L0Index ? L0Memory_56 : _GEN_61; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_63 = 6'h39 == L0Index ? L0Memory_57 : _GEN_62; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_64 = 6'h3a == L0Index ? L0Memory_58 : _GEN_63; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_65 = 6'h3b == L0Index ? L0Memory_59 : _GEN_64; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_66 = 6'h3c == L0Index ? L0Memory_60 : _GEN_65; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_67 = 6'h3d == L0Index ? L0Memory_61 : _GEN_66; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_68 = 6'h3e == L0Index ? L0Memory_62 : _GEN_67; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_69 = 6'h3f == L0Index ? L0Memory_63 : _GEN_68; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [6:0] _GEN_793 = {{1'd0}, L0Index}; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_70 = 7'h40 == _GEN_793 ? L0Memory_64 : _GEN_69; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_71 = 7'h41 == _GEN_793 ? L0Memory_65 : _GEN_70; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_72 = 7'h42 == _GEN_793 ? L0Memory_66 : _GEN_71; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_73 = 7'h43 == _GEN_793 ? L0Memory_67 : _GEN_72; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_74 = 7'h44 == _GEN_793 ? L0Memory_68 : _GEN_73; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_75 = 7'h45 == _GEN_793 ? L0Memory_69 : _GEN_74; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_76 = 7'h46 == _GEN_793 ? L0Memory_70 : _GEN_75; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_77 = 7'h47 == _GEN_793 ? L0Memory_71 : _GEN_76; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_78 = 7'h48 == _GEN_793 ? L0Memory_72 : _GEN_77; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_79 = 7'h49 == _GEN_793 ? L0Memory_73 : _GEN_78; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_80 = 7'h4a == _GEN_793 ? L0Memory_74 : _GEN_79; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_81 = 7'h4b == _GEN_793 ? L0Memory_75 : _GEN_80; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_82 = 7'h4c == _GEN_793 ? L0Memory_76 : _GEN_81; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_83 = 7'h4d == _GEN_793 ? L0Memory_77 : _GEN_82; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_84 = 7'h4e == _GEN_793 ? L0Memory_78 : _GEN_83; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_85 = 7'h4f == _GEN_793 ? L0Memory_79 : _GEN_84; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_86 = 7'h50 == _GEN_793 ? L0Memory_80 : _GEN_85; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_87 = 7'h51 == _GEN_793 ? L0Memory_81 : _GEN_86; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_88 = 7'h52 == _GEN_793 ? L0Memory_82 : _GEN_87; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_89 = 7'h53 == _GEN_793 ? L0Memory_83 : _GEN_88; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_90 = 7'h54 == _GEN_793 ? L0Memory_84 : _GEN_89; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_91 = 7'h55 == _GEN_793 ? L0Memory_85 : _GEN_90; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_92 = 7'h56 == _GEN_793 ? L0Memory_86 : _GEN_91; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_93 = 7'h57 == _GEN_793 ? L0Memory_87 : _GEN_92; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_94 = 7'h58 == _GEN_793 ? L0Memory_88 : _GEN_93; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_95 = 7'h59 == _GEN_793 ? L0Memory_89 : _GEN_94; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_96 = 7'h5a == _GEN_793 ? L0Memory_90 : _GEN_95; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_97 = 7'h5b == _GEN_793 ? L0Memory_91 : _GEN_96; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_98 = 7'h5c == _GEN_793 ? L0Memory_92 : _GEN_97; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_99 = 7'h5d == _GEN_793 ? L0Memory_93 : _GEN_98; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_100 = 7'h5e == _GEN_793 ? L0Memory_94 : _GEN_99; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_101 = 7'h5f == _GEN_793 ? L0Memory_95 : _GEN_100; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_102 = 7'h60 == _GEN_793 ? L0Memory_96 : _GEN_101; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_103 = 7'h61 == _GEN_793 ? L0Memory_97 : _GEN_102; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_104 = 7'h62 == _GEN_793 ? L0Memory_98 : _GEN_103; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_105 = 7'h63 == _GEN_793 ? L0Memory_99 : _GEN_104; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire  _GEN_575 = _T_12 ? 1'h0 : _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 157:12]
  wire  sel5 = _T_3 ? 1'h0 : _GEN_575; // @[Conditional.scala 40:58 PEArray.scala 112:12]
  reg [15:0] mux2out_reg; // @[PEArray.scala 90:28]
  reg [15:0] mux3out_reg; // @[PEArray.scala 91:28]
  reg [9:0] count; // @[PEArray.scala 101:22]
  reg [9:0] count_max; // @[PEArray.scala 102:22]
  reg [5:0] L0index_begin; // @[PEArray.scala 103:26]
  reg [5:0] GRU_out_width; // @[PEArray.scala 104:26]
  wire  _T_6 = 3'h0 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_7 = 3'h1 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_8 = 3'h2 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_9 = 3'h3 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_10 = 3'h4 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_11 = 3'h5 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_109 = _T_11 ? 3'h5 : state; // @[Conditional.scala 39:67 PEArray.scala 140:19 PEArray.scala 100:22]
  wire [2:0] _GEN_110 = _T_10 ? 3'h4 : _GEN_109; // @[Conditional.scala 39:67 PEArray.scala 136:19]
  wire [2:0] _GEN_111 = _T_9 ? 3'h3 : _GEN_110; // @[Conditional.scala 39:67 PEArray.scala 132:19]
  wire [2:0] _GEN_112 = _T_8 ? 3'h2 : _GEN_111; // @[Conditional.scala 39:67 PEArray.scala 128:19]
  wire [2:0] _GEN_113 = _T_7 ? 3'h1 : _GEN_112; // @[Conditional.scala 39:67 PEArray.scala 124:19]
  wire [7:0] _GEN_118 = io_control_signal_mask[6] ? io_control_signal_gru_out_width : {{2'd0}, GRU_out_width}; // @[PEArray.scala 116:57 PEArray.scala 145:23 PEArray.scala 104:26]
  wire [9:0] _count_T_1 = count + 10'h1; // @[PEArray.scala 162:24]
  wire [9:0] _GEN_120 = count != 10'h33 ? _count_T_1 : count; // @[PEArray.scala 161:27 PEArray.scala 162:15 PEArray.scala 101:22]
  wire [9:0] _GEN_124 = count != 10'h188 ? _count_T_1 : count; // @[PEArray.scala 183:28 PEArray.scala 184:15 PEArray.scala 101:22]
  wire [9:0] _GEN_125 = count == 10'h188 ? 10'h0 : _GEN_124; // @[PEArray.scala 186:28 PEArray.scala 187:15]
  wire [2:0] _GEN_126 = count == 10'h188 ? 3'h0 : state; // @[PEArray.scala 186:28 PEArray.scala 188:15 PEArray.scala 100:22]
  wire [9:0] _GEN_127 = count != count_max ? _count_T_1 : count; // @[PEArray.scala 192:32 PEArray.scala 193:15 PEArray.scala 101:22]
  wire [5:0] _GEN_128 = count == 10'h0 ? L0index_begin : L0Index; // @[PEArray.scala 195:26 PEArray.scala 196:17 PEArray.scala 39:24]
  wire [9:0] _T_27 = count_max - 10'h1; // @[PEArray.scala 198:51]
  wire [15:0] _GEN_129 = 6'h0 == L0Index ? io_FromL1 : L0Memory_0; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_130 = 6'h1 == L0Index ? io_FromL1 : L0Memory_1; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_131 = 6'h2 == L0Index ? io_FromL1 : L0Memory_2; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_132 = 6'h3 == L0Index ? io_FromL1 : L0Memory_3; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_133 = 6'h4 == L0Index ? io_FromL1 : L0Memory_4; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_134 = 6'h5 == L0Index ? io_FromL1 : L0Memory_5; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_135 = 6'h6 == L0Index ? io_FromL1 : L0Memory_6; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_136 = 6'h7 == L0Index ? io_FromL1 : L0Memory_7; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_137 = 6'h8 == L0Index ? io_FromL1 : L0Memory_8; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_138 = 6'h9 == L0Index ? io_FromL1 : L0Memory_9; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_139 = 6'ha == L0Index ? io_FromL1 : L0Memory_10; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_140 = 6'hb == L0Index ? io_FromL1 : L0Memory_11; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_141 = 6'hc == L0Index ? io_FromL1 : L0Memory_12; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_142 = 6'hd == L0Index ? io_FromL1 : L0Memory_13; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_143 = 6'he == L0Index ? io_FromL1 : L0Memory_14; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_144 = 6'hf == L0Index ? io_FromL1 : L0Memory_15; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_145 = 6'h10 == L0Index ? io_FromL1 : L0Memory_16; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_146 = 6'h11 == L0Index ? io_FromL1 : L0Memory_17; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_147 = 6'h12 == L0Index ? io_FromL1 : L0Memory_18; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_148 = 6'h13 == L0Index ? io_FromL1 : L0Memory_19; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_149 = 6'h14 == L0Index ? io_FromL1 : L0Memory_20; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_150 = 6'h15 == L0Index ? io_FromL1 : L0Memory_21; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_151 = 6'h16 == L0Index ? io_FromL1 : L0Memory_22; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_152 = 6'h17 == L0Index ? io_FromL1 : L0Memory_23; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_153 = 6'h18 == L0Index ? io_FromL1 : L0Memory_24; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_154 = 6'h19 == L0Index ? io_FromL1 : L0Memory_25; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_155 = 6'h1a == L0Index ? io_FromL1 : L0Memory_26; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_156 = 6'h1b == L0Index ? io_FromL1 : L0Memory_27; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_157 = 6'h1c == L0Index ? io_FromL1 : L0Memory_28; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_158 = 6'h1d == L0Index ? io_FromL1 : L0Memory_29; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_159 = 6'h1e == L0Index ? io_FromL1 : L0Memory_30; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_160 = 6'h1f == L0Index ? io_FromL1 : L0Memory_31; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_161 = 6'h20 == L0Index ? io_FromL1 : L0Memory_32; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_162 = 6'h21 == L0Index ? io_FromL1 : L0Memory_33; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_163 = 6'h22 == L0Index ? io_FromL1 : L0Memory_34; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_164 = 6'h23 == L0Index ? io_FromL1 : L0Memory_35; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_165 = 6'h24 == L0Index ? io_FromL1 : L0Memory_36; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_166 = 6'h25 == L0Index ? io_FromL1 : L0Memory_37; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_167 = 6'h26 == L0Index ? io_FromL1 : L0Memory_38; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_168 = 6'h27 == L0Index ? io_FromL1 : L0Memory_39; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_169 = 6'h28 == L0Index ? io_FromL1 : L0Memory_40; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_170 = 6'h29 == L0Index ? io_FromL1 : L0Memory_41; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_171 = 6'h2a == L0Index ? io_FromL1 : L0Memory_42; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_172 = 6'h2b == L0Index ? io_FromL1 : L0Memory_43; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_173 = 6'h2c == L0Index ? io_FromL1 : L0Memory_44; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_174 = 6'h2d == L0Index ? io_FromL1 : L0Memory_45; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_175 = 6'h2e == L0Index ? io_FromL1 : L0Memory_46; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_176 = 6'h2f == L0Index ? io_FromL1 : L0Memory_47; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_177 = 6'h30 == L0Index ? io_FromL1 : L0Memory_48; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_178 = 6'h31 == L0Index ? io_FromL1 : L0Memory_49; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_179 = 6'h32 == L0Index ? io_FromL1 : L0Memory_50; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_180 = 6'h33 == L0Index ? io_FromL1 : L0Memory_51; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_181 = 6'h34 == L0Index ? io_FromL1 : L0Memory_52; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_182 = 6'h35 == L0Index ? io_FromL1 : L0Memory_53; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_183 = 6'h36 == L0Index ? io_FromL1 : L0Memory_54; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_184 = 6'h37 == L0Index ? io_FromL1 : L0Memory_55; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_185 = 6'h38 == L0Index ? io_FromL1 : L0Memory_56; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_186 = 6'h39 == L0Index ? io_FromL1 : L0Memory_57; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_187 = 6'h3a == L0Index ? io_FromL1 : L0Memory_58; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_188 = 6'h3b == L0Index ? io_FromL1 : L0Memory_59; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_189 = 6'h3c == L0Index ? io_FromL1 : L0Memory_60; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_190 = 6'h3d == L0Index ? io_FromL1 : L0Memory_61; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_191 = 6'h3e == L0Index ? io_FromL1 : L0Memory_62; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_192 = 6'h3f == L0Index ? io_FromL1 : L0Memory_63; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_193 = 7'h40 == _GEN_793 ? io_FromL1 : L0Memory_64; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_194 = 7'h41 == _GEN_793 ? io_FromL1 : L0Memory_65; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_195 = 7'h42 == _GEN_793 ? io_FromL1 : L0Memory_66; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_196 = 7'h43 == _GEN_793 ? io_FromL1 : L0Memory_67; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_197 = 7'h44 == _GEN_793 ? io_FromL1 : L0Memory_68; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_198 = 7'h45 == _GEN_793 ? io_FromL1 : L0Memory_69; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_199 = 7'h46 == _GEN_793 ? io_FromL1 : L0Memory_70; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_200 = 7'h47 == _GEN_793 ? io_FromL1 : L0Memory_71; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_201 = 7'h48 == _GEN_793 ? io_FromL1 : L0Memory_72; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_202 = 7'h49 == _GEN_793 ? io_FromL1 : L0Memory_73; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_203 = 7'h4a == _GEN_793 ? io_FromL1 : L0Memory_74; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_204 = 7'h4b == _GEN_793 ? io_FromL1 : L0Memory_75; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_205 = 7'h4c == _GEN_793 ? io_FromL1 : L0Memory_76; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_206 = 7'h4d == _GEN_793 ? io_FromL1 : L0Memory_77; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_207 = 7'h4e == _GEN_793 ? io_FromL1 : L0Memory_78; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_208 = 7'h4f == _GEN_793 ? io_FromL1 : L0Memory_79; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_209 = 7'h50 == _GEN_793 ? io_FromL1 : L0Memory_80; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_210 = 7'h51 == _GEN_793 ? io_FromL1 : L0Memory_81; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_211 = 7'h52 == _GEN_793 ? io_FromL1 : L0Memory_82; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_212 = 7'h53 == _GEN_793 ? io_FromL1 : L0Memory_83; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_213 = 7'h54 == _GEN_793 ? io_FromL1 : L0Memory_84; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_214 = 7'h55 == _GEN_793 ? io_FromL1 : L0Memory_85; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_215 = 7'h56 == _GEN_793 ? io_FromL1 : L0Memory_86; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_216 = 7'h57 == _GEN_793 ? io_FromL1 : L0Memory_87; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_217 = 7'h58 == _GEN_793 ? io_FromL1 : L0Memory_88; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_218 = 7'h59 == _GEN_793 ? io_FromL1 : L0Memory_89; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_219 = 7'h5a == _GEN_793 ? io_FromL1 : L0Memory_90; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_220 = 7'h5b == _GEN_793 ? io_FromL1 : L0Memory_91; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_221 = 7'h5c == _GEN_793 ? io_FromL1 : L0Memory_92; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_222 = 7'h5d == _GEN_793 ? io_FromL1 : L0Memory_93; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_223 = 7'h5e == _GEN_793 ? io_FromL1 : L0Memory_94; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_224 = 7'h5f == _GEN_793 ? io_FromL1 : L0Memory_95; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_225 = 7'h60 == _GEN_793 ? io_FromL1 : L0Memory_96; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_226 = 7'h61 == _GEN_793 ? io_FromL1 : L0Memory_97; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_227 = 7'h62 == _GEN_793 ? io_FromL1 : L0Memory_98; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_228 = 7'h63 == _GEN_793 ? io_FromL1 : L0Memory_99; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [5:0] _L0Index_T_2 = L0Index + 6'h1; // @[PEArray.scala 200:28]
  wire [15:0] _GEN_229 = count >= 10'h1 & count <= _T_27 ? _GEN_129 : L0Memory_0; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_230 = count >= 10'h1 & count <= _T_27 ? _GEN_130 : L0Memory_1; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_231 = count >= 10'h1 & count <= _T_27 ? _GEN_131 : L0Memory_2; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_232 = count >= 10'h1 & count <= _T_27 ? _GEN_132 : L0Memory_3; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_233 = count >= 10'h1 & count <= _T_27 ? _GEN_133 : L0Memory_4; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_234 = count >= 10'h1 & count <= _T_27 ? _GEN_134 : L0Memory_5; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_235 = count >= 10'h1 & count <= _T_27 ? _GEN_135 : L0Memory_6; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_236 = count >= 10'h1 & count <= _T_27 ? _GEN_136 : L0Memory_7; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_237 = count >= 10'h1 & count <= _T_27 ? _GEN_137 : L0Memory_8; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_238 = count >= 10'h1 & count <= _T_27 ? _GEN_138 : L0Memory_9; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_239 = count >= 10'h1 & count <= _T_27 ? _GEN_139 : L0Memory_10; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_240 = count >= 10'h1 & count <= _T_27 ? _GEN_140 : L0Memory_11; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_241 = count >= 10'h1 & count <= _T_27 ? _GEN_141 : L0Memory_12; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_242 = count >= 10'h1 & count <= _T_27 ? _GEN_142 : L0Memory_13; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_243 = count >= 10'h1 & count <= _T_27 ? _GEN_143 : L0Memory_14; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_244 = count >= 10'h1 & count <= _T_27 ? _GEN_144 : L0Memory_15; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_245 = count >= 10'h1 & count <= _T_27 ? _GEN_145 : L0Memory_16; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_246 = count >= 10'h1 & count <= _T_27 ? _GEN_146 : L0Memory_17; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_247 = count >= 10'h1 & count <= _T_27 ? _GEN_147 : L0Memory_18; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_248 = count >= 10'h1 & count <= _T_27 ? _GEN_148 : L0Memory_19; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_249 = count >= 10'h1 & count <= _T_27 ? _GEN_149 : L0Memory_20; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_250 = count >= 10'h1 & count <= _T_27 ? _GEN_150 : L0Memory_21; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_251 = count >= 10'h1 & count <= _T_27 ? _GEN_151 : L0Memory_22; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_252 = count >= 10'h1 & count <= _T_27 ? _GEN_152 : L0Memory_23; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_253 = count >= 10'h1 & count <= _T_27 ? _GEN_153 : L0Memory_24; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_254 = count >= 10'h1 & count <= _T_27 ? _GEN_154 : L0Memory_25; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_255 = count >= 10'h1 & count <= _T_27 ? _GEN_155 : L0Memory_26; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_256 = count >= 10'h1 & count <= _T_27 ? _GEN_156 : L0Memory_27; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_257 = count >= 10'h1 & count <= _T_27 ? _GEN_157 : L0Memory_28; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_258 = count >= 10'h1 & count <= _T_27 ? _GEN_158 : L0Memory_29; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_259 = count >= 10'h1 & count <= _T_27 ? _GEN_159 : L0Memory_30; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_260 = count >= 10'h1 & count <= _T_27 ? _GEN_160 : L0Memory_31; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_261 = count >= 10'h1 & count <= _T_27 ? _GEN_161 : L0Memory_32; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_262 = count >= 10'h1 & count <= _T_27 ? _GEN_162 : L0Memory_33; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_263 = count >= 10'h1 & count <= _T_27 ? _GEN_163 : L0Memory_34; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_264 = count >= 10'h1 & count <= _T_27 ? _GEN_164 : L0Memory_35; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_265 = count >= 10'h1 & count <= _T_27 ? _GEN_165 : L0Memory_36; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_266 = count >= 10'h1 & count <= _T_27 ? _GEN_166 : L0Memory_37; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_267 = count >= 10'h1 & count <= _T_27 ? _GEN_167 : L0Memory_38; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_268 = count >= 10'h1 & count <= _T_27 ? _GEN_168 : L0Memory_39; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_269 = count >= 10'h1 & count <= _T_27 ? _GEN_169 : L0Memory_40; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_270 = count >= 10'h1 & count <= _T_27 ? _GEN_170 : L0Memory_41; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_271 = count >= 10'h1 & count <= _T_27 ? _GEN_171 : L0Memory_42; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_272 = count >= 10'h1 & count <= _T_27 ? _GEN_172 : L0Memory_43; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_273 = count >= 10'h1 & count <= _T_27 ? _GEN_173 : L0Memory_44; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_274 = count >= 10'h1 & count <= _T_27 ? _GEN_174 : L0Memory_45; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_275 = count >= 10'h1 & count <= _T_27 ? _GEN_175 : L0Memory_46; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_276 = count >= 10'h1 & count <= _T_27 ? _GEN_176 : L0Memory_47; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_277 = count >= 10'h1 & count <= _T_27 ? _GEN_177 : L0Memory_48; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_278 = count >= 10'h1 & count <= _T_27 ? _GEN_178 : L0Memory_49; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_279 = count >= 10'h1 & count <= _T_27 ? _GEN_179 : L0Memory_50; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_280 = count >= 10'h1 & count <= _T_27 ? _GEN_180 : L0Memory_51; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_281 = count >= 10'h1 & count <= _T_27 ? _GEN_181 : L0Memory_52; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_282 = count >= 10'h1 & count <= _T_27 ? _GEN_182 : L0Memory_53; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_283 = count >= 10'h1 & count <= _T_27 ? _GEN_183 : L0Memory_54; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_284 = count >= 10'h1 & count <= _T_27 ? _GEN_184 : L0Memory_55; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_285 = count >= 10'h1 & count <= _T_27 ? _GEN_185 : L0Memory_56; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_286 = count >= 10'h1 & count <= _T_27 ? _GEN_186 : L0Memory_57; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_287 = count >= 10'h1 & count <= _T_27 ? _GEN_187 : L0Memory_58; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_288 = count >= 10'h1 & count <= _T_27 ? _GEN_188 : L0Memory_59; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_289 = count >= 10'h1 & count <= _T_27 ? _GEN_189 : L0Memory_60; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_290 = count >= 10'h1 & count <= _T_27 ? _GEN_190 : L0Memory_61; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_291 = count >= 10'h1 & count <= _T_27 ? _GEN_191 : L0Memory_62; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_292 = count >= 10'h1 & count <= _T_27 ? _GEN_192 : L0Memory_63; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_293 = count >= 10'h1 & count <= _T_27 ? _GEN_193 : L0Memory_64; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_294 = count >= 10'h1 & count <= _T_27 ? _GEN_194 : L0Memory_65; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_295 = count >= 10'h1 & count <= _T_27 ? _GEN_195 : L0Memory_66; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_296 = count >= 10'h1 & count <= _T_27 ? _GEN_196 : L0Memory_67; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_297 = count >= 10'h1 & count <= _T_27 ? _GEN_197 : L0Memory_68; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_298 = count >= 10'h1 & count <= _T_27 ? _GEN_198 : L0Memory_69; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_299 = count >= 10'h1 & count <= _T_27 ? _GEN_199 : L0Memory_70; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_300 = count >= 10'h1 & count <= _T_27 ? _GEN_200 : L0Memory_71; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_301 = count >= 10'h1 & count <= _T_27 ? _GEN_201 : L0Memory_72; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_302 = count >= 10'h1 & count <= _T_27 ? _GEN_202 : L0Memory_73; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_303 = count >= 10'h1 & count <= _T_27 ? _GEN_203 : L0Memory_74; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_304 = count >= 10'h1 & count <= _T_27 ? _GEN_204 : L0Memory_75; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_305 = count >= 10'h1 & count <= _T_27 ? _GEN_205 : L0Memory_76; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_306 = count >= 10'h1 & count <= _T_27 ? _GEN_206 : L0Memory_77; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_307 = count >= 10'h1 & count <= _T_27 ? _GEN_207 : L0Memory_78; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_308 = count >= 10'h1 & count <= _T_27 ? _GEN_208 : L0Memory_79; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_309 = count >= 10'h1 & count <= _T_27 ? _GEN_209 : L0Memory_80; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_310 = count >= 10'h1 & count <= _T_27 ? _GEN_210 : L0Memory_81; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_311 = count >= 10'h1 & count <= _T_27 ? _GEN_211 : L0Memory_82; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_312 = count >= 10'h1 & count <= _T_27 ? _GEN_212 : L0Memory_83; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_313 = count >= 10'h1 & count <= _T_27 ? _GEN_213 : L0Memory_84; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_314 = count >= 10'h1 & count <= _T_27 ? _GEN_214 : L0Memory_85; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_315 = count >= 10'h1 & count <= _T_27 ? _GEN_215 : L0Memory_86; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_316 = count >= 10'h1 & count <= _T_27 ? _GEN_216 : L0Memory_87; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_317 = count >= 10'h1 & count <= _T_27 ? _GEN_217 : L0Memory_88; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_318 = count >= 10'h1 & count <= _T_27 ? _GEN_218 : L0Memory_89; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_319 = count >= 10'h1 & count <= _T_27 ? _GEN_219 : L0Memory_90; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_320 = count >= 10'h1 & count <= _T_27 ? _GEN_220 : L0Memory_91; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_321 = count >= 10'h1 & count <= _T_27 ? _GEN_221 : L0Memory_92; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_322 = count >= 10'h1 & count <= _T_27 ? _GEN_222 : L0Memory_93; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_323 = count >= 10'h1 & count <= _T_27 ? _GEN_223 : L0Memory_94; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_324 = count >= 10'h1 & count <= _T_27 ? _GEN_224 : L0Memory_95; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_325 = count >= 10'h1 & count <= _T_27 ? _GEN_225 : L0Memory_96; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_326 = count >= 10'h1 & count <= _T_27 ? _GEN_226 : L0Memory_97; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_327 = count >= 10'h1 & count <= _T_27 ? _GEN_227 : L0Memory_98; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_328 = count >= 10'h1 & count <= _T_27 ? _GEN_228 : L0Memory_99; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [5:0] _GEN_329 = count >= 10'h1 & count <= _T_27 ? _L0Index_T_2 : _GEN_128; // @[PEArray.scala 198:59 PEArray.scala 200:17]
  wire [9:0] _GEN_330 = count == count_max ? 10'h0 : _GEN_127; // @[PEArray.scala 202:32 PEArray.scala 203:15]
  wire [2:0] _GEN_331 = count == count_max ? 3'h0 : state; // @[PEArray.scala 202:32 PEArray.scala 204:15 PEArray.scala 100:22]
  wire [9:0] _GEN_865 = {{4'd0}, GRU_out_width}; // @[PEArray.scala 220:19]
  wire [9:0] _GEN_0 = count % _GEN_865; // @[PEArray.scala 220:19]
  wire [5:0] _T_36 = _GEN_0[5:0]; // @[PEArray.scala 220:19]
  wire [5:0] _T_38 = GRU_out_width - 6'h1; // @[PEArray.scala 220:55]
  wire [5:0] _GEN_334 = _T_36 == _T_38 ? _L0Index_T_2 : L0index_begin; // @[PEArray.scala 220:62 PEArray.scala 221:17 PEArray.scala 214:15]
  wire [5:0] _GEN_346 = _T_41 ? _GEN_334 : L0Index; // @[Conditional.scala 39:67 PEArray.scala 39:24]
  wire [9:0] _GEN_347 = _T_41 ? _GEN_330 : count; // @[Conditional.scala 39:67 PEArray.scala 101:22]
  wire [2:0] _GEN_348 = _T_41 ? _GEN_331 : state; // @[Conditional.scala 39:67 PEArray.scala 100:22]
  wire [5:0] _GEN_353 = _T_31 ? _GEN_334 : _GEN_346; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_354 = _T_31 ? _GEN_330 : _GEN_347; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_355 = _T_31 ? _GEN_331 : _GEN_348; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_356 = _T_22 ? _GEN_330 : _GEN_354; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_357 = _T_22 ? _GEN_329 : _GEN_353; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_458 = _T_22 ? _GEN_331 : _GEN_355; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_690 = _T_3 ? _GEN_118 : {{2'd0}, GRU_out_width}; // @[Conditional.scala 40:58 PEArray.scala 104:26]
  FP16MulAdder FP16MAC ( // @[PEArray.scala 72:23]
    .io_a(FP16MAC_io_a),
    .io_b(FP16MAC_io_b),
    .io_c(FP16MAC_io_c),
    .io_out(FP16MAC_io_out)
  );
  assign io_ToRightPE = mux3out_reg; // @[PEArray.scala 95:16]
  assign io_ToBelowPE = mux2out_reg; // @[PEArray.scala 94:16]
  assign FP16MAC_io_a = sel1 ? io_FromL1 : io_FromLeftPE; // @[PEArray.scala 50:14 PEArray.scala 50:23 PEArray.scala 51:24]
  assign FP16MAC_io_b = sel5 ? mux4out : _GEN_105; // @[PEArray.scala 77:13 PEArray.scala 78:18 PEArray.scala 81:18]
  assign FP16MAC_io_c = sel5 ? _GEN_105 : mux4out; // @[PEArray.scala 77:13 PEArray.scala 79:18 PEArray.scala 82:18]
  always @(posedge clock) begin
    if (reset) begin // @[PEArray.scala 39:24]
      L0Index <= 6'h0; // @[PEArray.scala 39:24]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h2; // @[PEArray.scala 159:15]
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h8; // @[PEArray.scala 181:15]
      end else begin
        L0Index <= _GEN_357;
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_0 <= _GEN_229;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_1 <= _GEN_230;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_2 <= _GEN_231;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_3 <= _GEN_232;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_4 <= _GEN_233;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_5 <= _GEN_234;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_6 <= _GEN_235;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_7 <= _GEN_236;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_8 <= _GEN_237;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_9 <= _GEN_238;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_10 <= _GEN_239;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_11 <= _GEN_240;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_12 <= _GEN_241;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_13 <= _GEN_242;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_14 <= _GEN_243;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_15 <= _GEN_244;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_16 <= _GEN_245;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_17 <= _GEN_246;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_18 <= _GEN_247;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_19 <= _GEN_248;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_20 <= _GEN_249;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_21 <= _GEN_250;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_22 <= _GEN_251;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_23 <= _GEN_252;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_24 <= _GEN_253;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_25 <= _GEN_254;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_26 <= _GEN_255;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_27 <= _GEN_256;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_28 <= _GEN_257;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_29 <= _GEN_258;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_30 <= _GEN_259;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_31 <= _GEN_260;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_32 <= _GEN_261;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_33 <= _GEN_262;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_34 <= _GEN_263;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_35 <= _GEN_264;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_36 <= _GEN_265;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_37 <= _GEN_266;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_38 <= _GEN_267;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_39 <= _GEN_268;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_40 <= _GEN_269;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_41 <= _GEN_270;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_42 <= _GEN_271;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_43 <= _GEN_272;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_44 <= _GEN_273;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_45 <= _GEN_274;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_46 <= _GEN_275;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_47 <= _GEN_276;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_48 <= _GEN_277;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_49 <= _GEN_278;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_50 <= _GEN_279;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_51 <= _GEN_280;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_52 <= _GEN_281;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_53 <= _GEN_282;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_54 <= _GEN_283;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_55 <= _GEN_284;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_56 <= _GEN_285;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_57 <= _GEN_286;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_58 <= _GEN_287;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_59 <= _GEN_288;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_60 <= _GEN_289;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_61 <= _GEN_290;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_62 <= _GEN_291;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_63 <= _GEN_292;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_64 <= _GEN_293;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_65 <= _GEN_294;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_66 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_67 <= _GEN_296;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_68 <= _GEN_297;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_69 <= _GEN_298;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_70 <= _GEN_299;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_71 <= _GEN_300;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_72 <= _GEN_301;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_73 <= _GEN_302;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_74 <= _GEN_303;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_75 <= _GEN_304;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_76 <= _GEN_305;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_77 <= _GEN_306;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_78 <= _GEN_307;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_79 <= _GEN_308;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_80 <= _GEN_309;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_81 <= _GEN_310;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_82 <= _GEN_311;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_83 <= _GEN_312;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_84 <= _GEN_313;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_85 <= _GEN_314;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_86 <= _GEN_315;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_87 <= _GEN_316;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_88 <= _GEN_317;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_89 <= _GEN_318;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_90 <= _GEN_319;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_91 <= _GEN_320;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_92 <= _GEN_321;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_93 <= _GEN_322;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_94 <= _GEN_323;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_95 <= _GEN_324;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_96 <= _GEN_325;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_97 <= _GEN_326;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_98 <= _GEN_327;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_99 <= _GEN_328;
          end
        end
      end
    end
    if (reset) begin // @[PEArray.scala 100:22]
      state <= 3'h0; // @[PEArray.scala 100:22]
    end else if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[6]) begin // @[PEArray.scala 116:57]
        if (_T_6) begin // @[Conditional.scala 40:58]
          state <= 3'h0; // @[PEArray.scala 120:19]
        end else begin
          state <= _GEN_113;
        end
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      if (count == 10'h33) begin // @[PEArray.scala 164:27]
        state <= 3'h0; // @[PEArray.scala 166:15]
      end
    end else if (_T_16) begin // @[Conditional.scala 39:67]
      state <= _GEN_126;
    end else begin
      state <= _GEN_458;
    end
    if (reset) begin // @[PEArray.scala 90:28]
      mux2out_reg <= 16'h0; // @[PEArray.scala 90:28]
    end else begin
      mux2out_reg <= MAC_out; // @[PEArray.scala 90:28]
    end
    if (reset) begin // @[PEArray.scala 91:28]
      mux3out_reg <= 16'h0; // @[PEArray.scala 91:28]
    end else if (sel3) begin // @[PEArray.scala 56:14]
      mux3out_reg <= MAC_out; // @[PEArray.scala 56:23]
    end else if (sel1) begin // @[PEArray.scala 50:14]
      mux3out_reg <= io_FromL1; // @[PEArray.scala 50:23]
    end else begin
      mux3out_reg <= io_FromLeftPE; // @[PEArray.scala 51:24]
    end
    if (reset) begin // @[PEArray.scala 101:22]
      count <= 10'h0; // @[PEArray.scala 101:22]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        if (count == 10'h33) begin // @[PEArray.scala 164:27]
          count <= 10'h0; // @[PEArray.scala 165:15]
        end else begin
          count <= _GEN_120;
        end
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        count <= _GEN_125;
      end else begin
        count <= _GEN_356;
      end
    end
    if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[6]) begin // @[PEArray.scala 116:57]
        count_max <= io_control_signal_count; // @[PEArray.scala 143:19]
      end
    end
    if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[6]) begin // @[PEArray.scala 116:57]
        L0index_begin <= io_control_signal_L0index; // @[PEArray.scala 144:23]
      end
    end
    GRU_out_width <= _GEN_690[5:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  L0Index = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  L0Memory_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  L0Memory_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  L0Memory_2 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  L0Memory_3 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  L0Memory_4 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  L0Memory_5 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  L0Memory_6 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  L0Memory_7 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  L0Memory_8 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  L0Memory_9 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  L0Memory_10 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  L0Memory_11 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  L0Memory_12 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  L0Memory_13 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  L0Memory_14 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  L0Memory_15 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  L0Memory_16 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  L0Memory_17 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  L0Memory_18 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  L0Memory_19 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  L0Memory_20 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  L0Memory_21 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  L0Memory_22 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  L0Memory_23 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  L0Memory_24 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  L0Memory_25 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  L0Memory_26 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  L0Memory_27 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  L0Memory_28 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  L0Memory_29 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  L0Memory_30 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  L0Memory_31 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  L0Memory_32 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  L0Memory_33 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  L0Memory_34 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  L0Memory_35 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  L0Memory_36 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  L0Memory_37 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  L0Memory_38 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  L0Memory_39 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  L0Memory_40 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  L0Memory_41 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  L0Memory_42 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  L0Memory_43 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  L0Memory_44 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  L0Memory_45 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  L0Memory_46 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  L0Memory_47 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  L0Memory_48 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  L0Memory_49 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  L0Memory_50 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  L0Memory_51 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  L0Memory_52 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  L0Memory_53 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  L0Memory_54 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  L0Memory_55 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  L0Memory_56 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  L0Memory_57 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  L0Memory_58 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  L0Memory_59 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  L0Memory_60 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  L0Memory_61 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  L0Memory_62 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  L0Memory_63 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  L0Memory_64 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  L0Memory_65 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  L0Memory_66 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  L0Memory_67 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  L0Memory_68 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  L0Memory_69 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  L0Memory_70 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  L0Memory_71 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  L0Memory_72 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  L0Memory_73 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  L0Memory_74 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  L0Memory_75 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  L0Memory_76 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  L0Memory_77 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  L0Memory_78 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  L0Memory_79 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  L0Memory_80 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  L0Memory_81 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  L0Memory_82 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  L0Memory_83 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  L0Memory_84 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  L0Memory_85 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  L0Memory_86 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  L0Memory_87 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  L0Memory_88 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  L0Memory_89 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  L0Memory_90 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  L0Memory_91 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  L0Memory_92 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  L0Memory_93 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  L0Memory_94 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  L0Memory_95 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  L0Memory_96 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  L0Memory_97 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  L0Memory_98 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  L0Memory_99 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  state = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  mux2out_reg = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  mux3out_reg = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  count = _RAND_104[9:0];
  _RAND_105 = {1{`RANDOM}};
  count_max = _RAND_105[9:0];
  _RAND_106 = {1{`RANDOM}};
  L0index_begin = _RAND_106[5:0];
  _RAND_107 = {1{`RANDOM}};
  GRU_out_width = _RAND_107[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PE_18(
  input         clock,
  input         reset,
  input  [15:0] io_FromAbovePE,
  input  [15:0] io_FromLeftPE,
  input  [15:0] io_FromL1,
  input  [11:0] io_control_signal_mask,
  output [15:0] io_ToRightPE,
  output [15:0] io_ToBelowPE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] FP16MAC_io_a; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_b; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_c; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_out; // @[PEArray.scala 72:23]
  reg [5:0] L0Index; // @[PEArray.scala 39:24]
  reg [15:0] L0Memory_0; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_1; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_2; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_3; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_4; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_5; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_6; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_7; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_8; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_9; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_10; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_11; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_12; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_13; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_14; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_15; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_16; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_17; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_18; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_19; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_20; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_21; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_22; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_23; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_24; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_25; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_26; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_27; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_28; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_29; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_30; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_31; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_32; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_33; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_34; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_35; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_36; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_37; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_38; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_39; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_40; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_41; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_42; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_43; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_44; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_45; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_46; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_47; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_48; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_49; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_50; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_51; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_52; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_53; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_54; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_55; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_56; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_57; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_58; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_59; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_60; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_61; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_62; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_63; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_64; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_65; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_66; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_67; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_68; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_69; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_70; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_71; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_72; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_73; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_74; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_75; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_76; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_77; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_78; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_79; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_80; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_81; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_82; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_83; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_84; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_85; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_86; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_87; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_88; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_89; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_90; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_91; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_92; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_93; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_94; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_95; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_96; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_97; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_98; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_99; // @[PEArray.scala 40:21]
  reg [2:0] state; // @[PEArray.scala 100:22]
  wire  _T_3 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_12 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_16 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_22 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_31 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_41 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_342 = _T_41 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 231:12 PEArray.scala 32:8]
  wire  _GEN_349 = _T_31 ? 1'h0 : _GEN_342; // @[Conditional.scala 39:67 PEArray.scala 208:12]
  wire  _GEN_459 = _T_22 | _GEN_349; // @[Conditional.scala 39:67 PEArray.scala 32:8]
  wire  _GEN_463 = _T_16 ? 1'h0 : _GEN_459; // @[Conditional.scala 39:67]
  wire  _GEN_572 = _T_12 | _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 149:12]
  wire  sel1 = _T_3 | _GEN_572; // @[Conditional.scala 40:58 PEArray.scala 108:12]
  wire [15:0] MAC_out = FP16MAC_io_out; // @[PEArray.scala 47:21 PEArray.scala 85:11]
  wire  _GEN_465 = _T_16 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 177:12]
  wire  _GEN_580 = _T_12 | _GEN_465; // @[Conditional.scala 39:67 PEArray.scala 34:8]
  wire  sel3 = _T_3 | _GEN_580; // @[Conditional.scala 40:58 PEArray.scala 110:12]
  wire [1:0] _GEN_344 = _T_41 ? 2'h2 : 2'h0; // @[Conditional.scala 39:67 PEArray.scala 233:12 PEArray.scala 35:8]
  wire [1:0] _GEN_351 = _T_31 ? 2'h2 : _GEN_344; // @[Conditional.scala 39:67 PEArray.scala 210:12]
  wire [1:0] _GEN_461 = _T_22 ? 2'h0 : _GEN_351; // @[Conditional.scala 39:67 PEArray.scala 35:8]
  wire [1:0] _GEN_466 = _T_16 ? 2'h0 : _GEN_461; // @[Conditional.scala 39:67 PEArray.scala 178:12]
  wire [1:0] _GEN_574 = _T_12 ? 2'h0 : _GEN_466; // @[Conditional.scala 39:67]
  wire [1:0] sel4 = _T_3 ? 2'h0 : _GEN_574; // @[Conditional.scala 40:58 PEArray.scala 111:12]
  wire [15:0] _GEN_3 = sel4 == 2'h2 ? io_FromL1 : 16'h0; // @[PEArray.scala 65:28 PEArray.scala 66:15 PEArray.scala 69:15]
  wire [15:0] _GEN_4 = sel4 == 2'h1 ? io_FromAbovePE : _GEN_3; // @[PEArray.scala 62:28 PEArray.scala 63:15]
  wire [15:0] mux4out = sel4 == 2'h0 ? 16'h0 : _GEN_4; // @[PEArray.scala 59:22 PEArray.scala 60:13]
  wire [15:0] _GEN_7 = 6'h1 == L0Index ? L0Memory_1 : L0Memory_0; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_8 = 6'h2 == L0Index ? L0Memory_2 : _GEN_7; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_9 = 6'h3 == L0Index ? L0Memory_3 : _GEN_8; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_10 = 6'h4 == L0Index ? L0Memory_4 : _GEN_9; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_11 = 6'h5 == L0Index ? L0Memory_5 : _GEN_10; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_12 = 6'h6 == L0Index ? L0Memory_6 : _GEN_11; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_13 = 6'h7 == L0Index ? L0Memory_7 : _GEN_12; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_14 = 6'h8 == L0Index ? L0Memory_8 : _GEN_13; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_15 = 6'h9 == L0Index ? L0Memory_9 : _GEN_14; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_16 = 6'ha == L0Index ? L0Memory_10 : _GEN_15; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_17 = 6'hb == L0Index ? L0Memory_11 : _GEN_16; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_18 = 6'hc == L0Index ? L0Memory_12 : _GEN_17; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_19 = 6'hd == L0Index ? L0Memory_13 : _GEN_18; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_20 = 6'he == L0Index ? L0Memory_14 : _GEN_19; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_21 = 6'hf == L0Index ? L0Memory_15 : _GEN_20; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_22 = 6'h10 == L0Index ? L0Memory_16 : _GEN_21; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_23 = 6'h11 == L0Index ? L0Memory_17 : _GEN_22; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_24 = 6'h12 == L0Index ? L0Memory_18 : _GEN_23; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_25 = 6'h13 == L0Index ? L0Memory_19 : _GEN_24; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_26 = 6'h14 == L0Index ? L0Memory_20 : _GEN_25; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_27 = 6'h15 == L0Index ? L0Memory_21 : _GEN_26; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_28 = 6'h16 == L0Index ? L0Memory_22 : _GEN_27; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_29 = 6'h17 == L0Index ? L0Memory_23 : _GEN_28; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_30 = 6'h18 == L0Index ? L0Memory_24 : _GEN_29; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_31 = 6'h19 == L0Index ? L0Memory_25 : _GEN_30; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_32 = 6'h1a == L0Index ? L0Memory_26 : _GEN_31; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_33 = 6'h1b == L0Index ? L0Memory_27 : _GEN_32; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_34 = 6'h1c == L0Index ? L0Memory_28 : _GEN_33; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_35 = 6'h1d == L0Index ? L0Memory_29 : _GEN_34; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_36 = 6'h1e == L0Index ? L0Memory_30 : _GEN_35; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_37 = 6'h1f == L0Index ? L0Memory_31 : _GEN_36; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_38 = 6'h20 == L0Index ? L0Memory_32 : _GEN_37; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_39 = 6'h21 == L0Index ? L0Memory_33 : _GEN_38; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_40 = 6'h22 == L0Index ? L0Memory_34 : _GEN_39; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_41 = 6'h23 == L0Index ? L0Memory_35 : _GEN_40; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_42 = 6'h24 == L0Index ? L0Memory_36 : _GEN_41; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_43 = 6'h25 == L0Index ? L0Memory_37 : _GEN_42; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_44 = 6'h26 == L0Index ? L0Memory_38 : _GEN_43; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_45 = 6'h27 == L0Index ? L0Memory_39 : _GEN_44; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_46 = 6'h28 == L0Index ? L0Memory_40 : _GEN_45; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_47 = 6'h29 == L0Index ? L0Memory_41 : _GEN_46; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_48 = 6'h2a == L0Index ? L0Memory_42 : _GEN_47; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_49 = 6'h2b == L0Index ? L0Memory_43 : _GEN_48; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_50 = 6'h2c == L0Index ? L0Memory_44 : _GEN_49; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_51 = 6'h2d == L0Index ? L0Memory_45 : _GEN_50; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_52 = 6'h2e == L0Index ? L0Memory_46 : _GEN_51; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_53 = 6'h2f == L0Index ? L0Memory_47 : _GEN_52; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_54 = 6'h30 == L0Index ? L0Memory_48 : _GEN_53; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_55 = 6'h31 == L0Index ? L0Memory_49 : _GEN_54; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_56 = 6'h32 == L0Index ? L0Memory_50 : _GEN_55; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_57 = 6'h33 == L0Index ? L0Memory_51 : _GEN_56; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_58 = 6'h34 == L0Index ? L0Memory_52 : _GEN_57; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_59 = 6'h35 == L0Index ? L0Memory_53 : _GEN_58; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_60 = 6'h36 == L0Index ? L0Memory_54 : _GEN_59; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_61 = 6'h37 == L0Index ? L0Memory_55 : _GEN_60; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_62 = 6'h38 == L0Index ? L0Memory_56 : _GEN_61; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_63 = 6'h39 == L0Index ? L0Memory_57 : _GEN_62; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_64 = 6'h3a == L0Index ? L0Memory_58 : _GEN_63; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_65 = 6'h3b == L0Index ? L0Memory_59 : _GEN_64; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_66 = 6'h3c == L0Index ? L0Memory_60 : _GEN_65; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_67 = 6'h3d == L0Index ? L0Memory_61 : _GEN_66; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_68 = 6'h3e == L0Index ? L0Memory_62 : _GEN_67; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_69 = 6'h3f == L0Index ? L0Memory_63 : _GEN_68; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [6:0] _GEN_793 = {{1'd0}, L0Index}; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_70 = 7'h40 == _GEN_793 ? L0Memory_64 : _GEN_69; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_71 = 7'h41 == _GEN_793 ? L0Memory_65 : _GEN_70; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_72 = 7'h42 == _GEN_793 ? L0Memory_66 : _GEN_71; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_73 = 7'h43 == _GEN_793 ? L0Memory_67 : _GEN_72; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_74 = 7'h44 == _GEN_793 ? L0Memory_68 : _GEN_73; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_75 = 7'h45 == _GEN_793 ? L0Memory_69 : _GEN_74; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_76 = 7'h46 == _GEN_793 ? L0Memory_70 : _GEN_75; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_77 = 7'h47 == _GEN_793 ? L0Memory_71 : _GEN_76; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_78 = 7'h48 == _GEN_793 ? L0Memory_72 : _GEN_77; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_79 = 7'h49 == _GEN_793 ? L0Memory_73 : _GEN_78; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_80 = 7'h4a == _GEN_793 ? L0Memory_74 : _GEN_79; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_81 = 7'h4b == _GEN_793 ? L0Memory_75 : _GEN_80; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_82 = 7'h4c == _GEN_793 ? L0Memory_76 : _GEN_81; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_83 = 7'h4d == _GEN_793 ? L0Memory_77 : _GEN_82; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_84 = 7'h4e == _GEN_793 ? L0Memory_78 : _GEN_83; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_85 = 7'h4f == _GEN_793 ? L0Memory_79 : _GEN_84; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_86 = 7'h50 == _GEN_793 ? L0Memory_80 : _GEN_85; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_87 = 7'h51 == _GEN_793 ? L0Memory_81 : _GEN_86; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_88 = 7'h52 == _GEN_793 ? L0Memory_82 : _GEN_87; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_89 = 7'h53 == _GEN_793 ? L0Memory_83 : _GEN_88; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_90 = 7'h54 == _GEN_793 ? L0Memory_84 : _GEN_89; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_91 = 7'h55 == _GEN_793 ? L0Memory_85 : _GEN_90; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_92 = 7'h56 == _GEN_793 ? L0Memory_86 : _GEN_91; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_93 = 7'h57 == _GEN_793 ? L0Memory_87 : _GEN_92; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_94 = 7'h58 == _GEN_793 ? L0Memory_88 : _GEN_93; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_95 = 7'h59 == _GEN_793 ? L0Memory_89 : _GEN_94; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_96 = 7'h5a == _GEN_793 ? L0Memory_90 : _GEN_95; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_97 = 7'h5b == _GEN_793 ? L0Memory_91 : _GEN_96; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_98 = 7'h5c == _GEN_793 ? L0Memory_92 : _GEN_97; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_99 = 7'h5d == _GEN_793 ? L0Memory_93 : _GEN_98; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_100 = 7'h5e == _GEN_793 ? L0Memory_94 : _GEN_99; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_101 = 7'h5f == _GEN_793 ? L0Memory_95 : _GEN_100; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_102 = 7'h60 == _GEN_793 ? L0Memory_96 : _GEN_101; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_103 = 7'h61 == _GEN_793 ? L0Memory_97 : _GEN_102; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_104 = 7'h62 == _GEN_793 ? L0Memory_98 : _GEN_103; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_105 = 7'h63 == _GEN_793 ? L0Memory_99 : _GEN_104; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire  _GEN_575 = _T_12 ? 1'h0 : _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 157:12]
  wire  sel5 = _T_3 ? 1'h0 : _GEN_575; // @[Conditional.scala 40:58 PEArray.scala 112:12]
  reg [15:0] mux2out_reg; // @[PEArray.scala 90:28]
  reg [15:0] mux3out_reg; // @[PEArray.scala 91:28]
  reg [9:0] count; // @[PEArray.scala 101:22]
  reg [5:0] GRU_out_width; // @[PEArray.scala 104:26]
  wire [7:0] _GEN_118 = io_control_signal_mask[5] ? 8'h0 : {{2'd0}, GRU_out_width}; // @[PEArray.scala 116:57 PEArray.scala 145:23 PEArray.scala 104:26]
  wire [9:0] _count_T_1 = count + 10'h1; // @[PEArray.scala 162:24]
  wire [9:0] _GEN_120 = count != 10'h33 ? _count_T_1 : count; // @[PEArray.scala 161:27 PEArray.scala 162:15 PEArray.scala 101:22]
  wire [9:0] _GEN_124 = count != 10'h188 ? _count_T_1 : count; // @[PEArray.scala 183:28 PEArray.scala 184:15 PEArray.scala 101:22]
  wire [9:0] _GEN_125 = count == 10'h188 ? 10'h0 : _GEN_124; // @[PEArray.scala 186:28 PEArray.scala 187:15]
  wire [2:0] _GEN_126 = count == 10'h188 ? 3'h0 : state; // @[PEArray.scala 186:28 PEArray.scala 188:15 PEArray.scala 100:22]
  wire [9:0] _GEN_127 = count != 10'h0 ? _count_T_1 : count; // @[PEArray.scala 192:32 PEArray.scala 193:15 PEArray.scala 101:22]
  wire  _T_24 = count == 10'h0; // @[PEArray.scala 195:18]
  wire [5:0] _GEN_128 = count == 10'h0 ? 6'h0 : L0Index; // @[PEArray.scala 195:26 PEArray.scala 196:17 PEArray.scala 39:24]
  wire [9:0] _T_27 = 10'h0 - 10'h1; // @[PEArray.scala 198:51]
  wire [15:0] _GEN_129 = 6'h0 == L0Index ? io_FromL1 : L0Memory_0; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_130 = 6'h1 == L0Index ? io_FromL1 : L0Memory_1; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_131 = 6'h2 == L0Index ? io_FromL1 : L0Memory_2; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_132 = 6'h3 == L0Index ? io_FromL1 : L0Memory_3; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_133 = 6'h4 == L0Index ? io_FromL1 : L0Memory_4; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_134 = 6'h5 == L0Index ? io_FromL1 : L0Memory_5; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_135 = 6'h6 == L0Index ? io_FromL1 : L0Memory_6; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_136 = 6'h7 == L0Index ? io_FromL1 : L0Memory_7; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_137 = 6'h8 == L0Index ? io_FromL1 : L0Memory_8; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_138 = 6'h9 == L0Index ? io_FromL1 : L0Memory_9; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_139 = 6'ha == L0Index ? io_FromL1 : L0Memory_10; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_140 = 6'hb == L0Index ? io_FromL1 : L0Memory_11; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_141 = 6'hc == L0Index ? io_FromL1 : L0Memory_12; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_142 = 6'hd == L0Index ? io_FromL1 : L0Memory_13; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_143 = 6'he == L0Index ? io_FromL1 : L0Memory_14; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_144 = 6'hf == L0Index ? io_FromL1 : L0Memory_15; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_145 = 6'h10 == L0Index ? io_FromL1 : L0Memory_16; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_146 = 6'h11 == L0Index ? io_FromL1 : L0Memory_17; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_147 = 6'h12 == L0Index ? io_FromL1 : L0Memory_18; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_148 = 6'h13 == L0Index ? io_FromL1 : L0Memory_19; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_149 = 6'h14 == L0Index ? io_FromL1 : L0Memory_20; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_150 = 6'h15 == L0Index ? io_FromL1 : L0Memory_21; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_151 = 6'h16 == L0Index ? io_FromL1 : L0Memory_22; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_152 = 6'h17 == L0Index ? io_FromL1 : L0Memory_23; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_153 = 6'h18 == L0Index ? io_FromL1 : L0Memory_24; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_154 = 6'h19 == L0Index ? io_FromL1 : L0Memory_25; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_155 = 6'h1a == L0Index ? io_FromL1 : L0Memory_26; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_156 = 6'h1b == L0Index ? io_FromL1 : L0Memory_27; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_157 = 6'h1c == L0Index ? io_FromL1 : L0Memory_28; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_158 = 6'h1d == L0Index ? io_FromL1 : L0Memory_29; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_159 = 6'h1e == L0Index ? io_FromL1 : L0Memory_30; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_160 = 6'h1f == L0Index ? io_FromL1 : L0Memory_31; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_161 = 6'h20 == L0Index ? io_FromL1 : L0Memory_32; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_162 = 6'h21 == L0Index ? io_FromL1 : L0Memory_33; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_163 = 6'h22 == L0Index ? io_FromL1 : L0Memory_34; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_164 = 6'h23 == L0Index ? io_FromL1 : L0Memory_35; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_165 = 6'h24 == L0Index ? io_FromL1 : L0Memory_36; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_166 = 6'h25 == L0Index ? io_FromL1 : L0Memory_37; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_167 = 6'h26 == L0Index ? io_FromL1 : L0Memory_38; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_168 = 6'h27 == L0Index ? io_FromL1 : L0Memory_39; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_169 = 6'h28 == L0Index ? io_FromL1 : L0Memory_40; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_170 = 6'h29 == L0Index ? io_FromL1 : L0Memory_41; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_171 = 6'h2a == L0Index ? io_FromL1 : L0Memory_42; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_172 = 6'h2b == L0Index ? io_FromL1 : L0Memory_43; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_173 = 6'h2c == L0Index ? io_FromL1 : L0Memory_44; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_174 = 6'h2d == L0Index ? io_FromL1 : L0Memory_45; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_175 = 6'h2e == L0Index ? io_FromL1 : L0Memory_46; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_176 = 6'h2f == L0Index ? io_FromL1 : L0Memory_47; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_177 = 6'h30 == L0Index ? io_FromL1 : L0Memory_48; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_178 = 6'h31 == L0Index ? io_FromL1 : L0Memory_49; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_179 = 6'h32 == L0Index ? io_FromL1 : L0Memory_50; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_180 = 6'h33 == L0Index ? io_FromL1 : L0Memory_51; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_181 = 6'h34 == L0Index ? io_FromL1 : L0Memory_52; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_182 = 6'h35 == L0Index ? io_FromL1 : L0Memory_53; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_183 = 6'h36 == L0Index ? io_FromL1 : L0Memory_54; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_184 = 6'h37 == L0Index ? io_FromL1 : L0Memory_55; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_185 = 6'h38 == L0Index ? io_FromL1 : L0Memory_56; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_186 = 6'h39 == L0Index ? io_FromL1 : L0Memory_57; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_187 = 6'h3a == L0Index ? io_FromL1 : L0Memory_58; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_188 = 6'h3b == L0Index ? io_FromL1 : L0Memory_59; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_189 = 6'h3c == L0Index ? io_FromL1 : L0Memory_60; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_190 = 6'h3d == L0Index ? io_FromL1 : L0Memory_61; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_191 = 6'h3e == L0Index ? io_FromL1 : L0Memory_62; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_192 = 6'h3f == L0Index ? io_FromL1 : L0Memory_63; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_193 = 7'h40 == _GEN_793 ? io_FromL1 : L0Memory_64; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_194 = 7'h41 == _GEN_793 ? io_FromL1 : L0Memory_65; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_195 = 7'h42 == _GEN_793 ? io_FromL1 : L0Memory_66; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_196 = 7'h43 == _GEN_793 ? io_FromL1 : L0Memory_67; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_197 = 7'h44 == _GEN_793 ? io_FromL1 : L0Memory_68; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_198 = 7'h45 == _GEN_793 ? io_FromL1 : L0Memory_69; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_199 = 7'h46 == _GEN_793 ? io_FromL1 : L0Memory_70; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_200 = 7'h47 == _GEN_793 ? io_FromL1 : L0Memory_71; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_201 = 7'h48 == _GEN_793 ? io_FromL1 : L0Memory_72; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_202 = 7'h49 == _GEN_793 ? io_FromL1 : L0Memory_73; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_203 = 7'h4a == _GEN_793 ? io_FromL1 : L0Memory_74; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_204 = 7'h4b == _GEN_793 ? io_FromL1 : L0Memory_75; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_205 = 7'h4c == _GEN_793 ? io_FromL1 : L0Memory_76; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_206 = 7'h4d == _GEN_793 ? io_FromL1 : L0Memory_77; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_207 = 7'h4e == _GEN_793 ? io_FromL1 : L0Memory_78; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_208 = 7'h4f == _GEN_793 ? io_FromL1 : L0Memory_79; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_209 = 7'h50 == _GEN_793 ? io_FromL1 : L0Memory_80; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_210 = 7'h51 == _GEN_793 ? io_FromL1 : L0Memory_81; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_211 = 7'h52 == _GEN_793 ? io_FromL1 : L0Memory_82; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_212 = 7'h53 == _GEN_793 ? io_FromL1 : L0Memory_83; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_213 = 7'h54 == _GEN_793 ? io_FromL1 : L0Memory_84; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_214 = 7'h55 == _GEN_793 ? io_FromL1 : L0Memory_85; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_215 = 7'h56 == _GEN_793 ? io_FromL1 : L0Memory_86; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_216 = 7'h57 == _GEN_793 ? io_FromL1 : L0Memory_87; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_217 = 7'h58 == _GEN_793 ? io_FromL1 : L0Memory_88; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_218 = 7'h59 == _GEN_793 ? io_FromL1 : L0Memory_89; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_219 = 7'h5a == _GEN_793 ? io_FromL1 : L0Memory_90; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_220 = 7'h5b == _GEN_793 ? io_FromL1 : L0Memory_91; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_221 = 7'h5c == _GEN_793 ? io_FromL1 : L0Memory_92; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_222 = 7'h5d == _GEN_793 ? io_FromL1 : L0Memory_93; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_223 = 7'h5e == _GEN_793 ? io_FromL1 : L0Memory_94; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_224 = 7'h5f == _GEN_793 ? io_FromL1 : L0Memory_95; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_225 = 7'h60 == _GEN_793 ? io_FromL1 : L0Memory_96; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_226 = 7'h61 == _GEN_793 ? io_FromL1 : L0Memory_97; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_227 = 7'h62 == _GEN_793 ? io_FromL1 : L0Memory_98; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_228 = 7'h63 == _GEN_793 ? io_FromL1 : L0Memory_99; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [5:0] _L0Index_T_2 = L0Index + 6'h1; // @[PEArray.scala 200:28]
  wire [15:0] _GEN_229 = count >= 10'h1 & count <= _T_27 ? _GEN_129 : L0Memory_0; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_230 = count >= 10'h1 & count <= _T_27 ? _GEN_130 : L0Memory_1; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_231 = count >= 10'h1 & count <= _T_27 ? _GEN_131 : L0Memory_2; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_232 = count >= 10'h1 & count <= _T_27 ? _GEN_132 : L0Memory_3; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_233 = count >= 10'h1 & count <= _T_27 ? _GEN_133 : L0Memory_4; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_234 = count >= 10'h1 & count <= _T_27 ? _GEN_134 : L0Memory_5; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_235 = count >= 10'h1 & count <= _T_27 ? _GEN_135 : L0Memory_6; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_236 = count >= 10'h1 & count <= _T_27 ? _GEN_136 : L0Memory_7; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_237 = count >= 10'h1 & count <= _T_27 ? _GEN_137 : L0Memory_8; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_238 = count >= 10'h1 & count <= _T_27 ? _GEN_138 : L0Memory_9; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_239 = count >= 10'h1 & count <= _T_27 ? _GEN_139 : L0Memory_10; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_240 = count >= 10'h1 & count <= _T_27 ? _GEN_140 : L0Memory_11; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_241 = count >= 10'h1 & count <= _T_27 ? _GEN_141 : L0Memory_12; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_242 = count >= 10'h1 & count <= _T_27 ? _GEN_142 : L0Memory_13; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_243 = count >= 10'h1 & count <= _T_27 ? _GEN_143 : L0Memory_14; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_244 = count >= 10'h1 & count <= _T_27 ? _GEN_144 : L0Memory_15; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_245 = count >= 10'h1 & count <= _T_27 ? _GEN_145 : L0Memory_16; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_246 = count >= 10'h1 & count <= _T_27 ? _GEN_146 : L0Memory_17; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_247 = count >= 10'h1 & count <= _T_27 ? _GEN_147 : L0Memory_18; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_248 = count >= 10'h1 & count <= _T_27 ? _GEN_148 : L0Memory_19; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_249 = count >= 10'h1 & count <= _T_27 ? _GEN_149 : L0Memory_20; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_250 = count >= 10'h1 & count <= _T_27 ? _GEN_150 : L0Memory_21; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_251 = count >= 10'h1 & count <= _T_27 ? _GEN_151 : L0Memory_22; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_252 = count >= 10'h1 & count <= _T_27 ? _GEN_152 : L0Memory_23; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_253 = count >= 10'h1 & count <= _T_27 ? _GEN_153 : L0Memory_24; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_254 = count >= 10'h1 & count <= _T_27 ? _GEN_154 : L0Memory_25; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_255 = count >= 10'h1 & count <= _T_27 ? _GEN_155 : L0Memory_26; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_256 = count >= 10'h1 & count <= _T_27 ? _GEN_156 : L0Memory_27; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_257 = count >= 10'h1 & count <= _T_27 ? _GEN_157 : L0Memory_28; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_258 = count >= 10'h1 & count <= _T_27 ? _GEN_158 : L0Memory_29; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_259 = count >= 10'h1 & count <= _T_27 ? _GEN_159 : L0Memory_30; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_260 = count >= 10'h1 & count <= _T_27 ? _GEN_160 : L0Memory_31; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_261 = count >= 10'h1 & count <= _T_27 ? _GEN_161 : L0Memory_32; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_262 = count >= 10'h1 & count <= _T_27 ? _GEN_162 : L0Memory_33; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_263 = count >= 10'h1 & count <= _T_27 ? _GEN_163 : L0Memory_34; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_264 = count >= 10'h1 & count <= _T_27 ? _GEN_164 : L0Memory_35; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_265 = count >= 10'h1 & count <= _T_27 ? _GEN_165 : L0Memory_36; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_266 = count >= 10'h1 & count <= _T_27 ? _GEN_166 : L0Memory_37; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_267 = count >= 10'h1 & count <= _T_27 ? _GEN_167 : L0Memory_38; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_268 = count >= 10'h1 & count <= _T_27 ? _GEN_168 : L0Memory_39; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_269 = count >= 10'h1 & count <= _T_27 ? _GEN_169 : L0Memory_40; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_270 = count >= 10'h1 & count <= _T_27 ? _GEN_170 : L0Memory_41; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_271 = count >= 10'h1 & count <= _T_27 ? _GEN_171 : L0Memory_42; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_272 = count >= 10'h1 & count <= _T_27 ? _GEN_172 : L0Memory_43; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_273 = count >= 10'h1 & count <= _T_27 ? _GEN_173 : L0Memory_44; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_274 = count >= 10'h1 & count <= _T_27 ? _GEN_174 : L0Memory_45; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_275 = count >= 10'h1 & count <= _T_27 ? _GEN_175 : L0Memory_46; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_276 = count >= 10'h1 & count <= _T_27 ? _GEN_176 : L0Memory_47; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_277 = count >= 10'h1 & count <= _T_27 ? _GEN_177 : L0Memory_48; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_278 = count >= 10'h1 & count <= _T_27 ? _GEN_178 : L0Memory_49; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_279 = count >= 10'h1 & count <= _T_27 ? _GEN_179 : L0Memory_50; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_280 = count >= 10'h1 & count <= _T_27 ? _GEN_180 : L0Memory_51; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_281 = count >= 10'h1 & count <= _T_27 ? _GEN_181 : L0Memory_52; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_282 = count >= 10'h1 & count <= _T_27 ? _GEN_182 : L0Memory_53; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_283 = count >= 10'h1 & count <= _T_27 ? _GEN_183 : L0Memory_54; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_284 = count >= 10'h1 & count <= _T_27 ? _GEN_184 : L0Memory_55; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_285 = count >= 10'h1 & count <= _T_27 ? _GEN_185 : L0Memory_56; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_286 = count >= 10'h1 & count <= _T_27 ? _GEN_186 : L0Memory_57; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_287 = count >= 10'h1 & count <= _T_27 ? _GEN_187 : L0Memory_58; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_288 = count >= 10'h1 & count <= _T_27 ? _GEN_188 : L0Memory_59; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_289 = count >= 10'h1 & count <= _T_27 ? _GEN_189 : L0Memory_60; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_290 = count >= 10'h1 & count <= _T_27 ? _GEN_190 : L0Memory_61; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_291 = count >= 10'h1 & count <= _T_27 ? _GEN_191 : L0Memory_62; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_292 = count >= 10'h1 & count <= _T_27 ? _GEN_192 : L0Memory_63; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_293 = count >= 10'h1 & count <= _T_27 ? _GEN_193 : L0Memory_64; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_294 = count >= 10'h1 & count <= _T_27 ? _GEN_194 : L0Memory_65; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_295 = count >= 10'h1 & count <= _T_27 ? _GEN_195 : L0Memory_66; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_296 = count >= 10'h1 & count <= _T_27 ? _GEN_196 : L0Memory_67; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_297 = count >= 10'h1 & count <= _T_27 ? _GEN_197 : L0Memory_68; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_298 = count >= 10'h1 & count <= _T_27 ? _GEN_198 : L0Memory_69; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_299 = count >= 10'h1 & count <= _T_27 ? _GEN_199 : L0Memory_70; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_300 = count >= 10'h1 & count <= _T_27 ? _GEN_200 : L0Memory_71; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_301 = count >= 10'h1 & count <= _T_27 ? _GEN_201 : L0Memory_72; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_302 = count >= 10'h1 & count <= _T_27 ? _GEN_202 : L0Memory_73; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_303 = count >= 10'h1 & count <= _T_27 ? _GEN_203 : L0Memory_74; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_304 = count >= 10'h1 & count <= _T_27 ? _GEN_204 : L0Memory_75; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_305 = count >= 10'h1 & count <= _T_27 ? _GEN_205 : L0Memory_76; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_306 = count >= 10'h1 & count <= _T_27 ? _GEN_206 : L0Memory_77; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_307 = count >= 10'h1 & count <= _T_27 ? _GEN_207 : L0Memory_78; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_308 = count >= 10'h1 & count <= _T_27 ? _GEN_208 : L0Memory_79; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_309 = count >= 10'h1 & count <= _T_27 ? _GEN_209 : L0Memory_80; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_310 = count >= 10'h1 & count <= _T_27 ? _GEN_210 : L0Memory_81; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_311 = count >= 10'h1 & count <= _T_27 ? _GEN_211 : L0Memory_82; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_312 = count >= 10'h1 & count <= _T_27 ? _GEN_212 : L0Memory_83; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_313 = count >= 10'h1 & count <= _T_27 ? _GEN_213 : L0Memory_84; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_314 = count >= 10'h1 & count <= _T_27 ? _GEN_214 : L0Memory_85; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_315 = count >= 10'h1 & count <= _T_27 ? _GEN_215 : L0Memory_86; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_316 = count >= 10'h1 & count <= _T_27 ? _GEN_216 : L0Memory_87; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_317 = count >= 10'h1 & count <= _T_27 ? _GEN_217 : L0Memory_88; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_318 = count >= 10'h1 & count <= _T_27 ? _GEN_218 : L0Memory_89; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_319 = count >= 10'h1 & count <= _T_27 ? _GEN_219 : L0Memory_90; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_320 = count >= 10'h1 & count <= _T_27 ? _GEN_220 : L0Memory_91; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_321 = count >= 10'h1 & count <= _T_27 ? _GEN_221 : L0Memory_92; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_322 = count >= 10'h1 & count <= _T_27 ? _GEN_222 : L0Memory_93; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_323 = count >= 10'h1 & count <= _T_27 ? _GEN_223 : L0Memory_94; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_324 = count >= 10'h1 & count <= _T_27 ? _GEN_224 : L0Memory_95; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_325 = count >= 10'h1 & count <= _T_27 ? _GEN_225 : L0Memory_96; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_326 = count >= 10'h1 & count <= _T_27 ? _GEN_226 : L0Memory_97; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_327 = count >= 10'h1 & count <= _T_27 ? _GEN_227 : L0Memory_98; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_328 = count >= 10'h1 & count <= _T_27 ? _GEN_228 : L0Memory_99; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [5:0] _GEN_329 = count >= 10'h1 & count <= _T_27 ? _L0Index_T_2 : _GEN_128; // @[PEArray.scala 198:59 PEArray.scala 200:17]
  wire [9:0] _GEN_330 = _T_24 ? 10'h0 : _GEN_127; // @[PEArray.scala 202:32 PEArray.scala 203:15]
  wire [2:0] _GEN_331 = _T_24 ? 3'h0 : state; // @[PEArray.scala 202:32 PEArray.scala 204:15 PEArray.scala 100:22]
  wire [9:0] _GEN_865 = {{4'd0}, GRU_out_width}; // @[PEArray.scala 220:19]
  wire [9:0] _GEN_0 = count % _GEN_865; // @[PEArray.scala 220:19]
  wire [5:0] _T_36 = _GEN_0[5:0]; // @[PEArray.scala 220:19]
  wire [5:0] _T_38 = GRU_out_width - 6'h1; // @[PEArray.scala 220:55]
  wire [5:0] _GEN_334 = _T_36 == _T_38 ? _L0Index_T_2 : 6'h0; // @[PEArray.scala 220:62 PEArray.scala 221:17 PEArray.scala 214:15]
  wire [5:0] _GEN_346 = _T_41 ? _GEN_334 : L0Index; // @[Conditional.scala 39:67 PEArray.scala 39:24]
  wire [9:0] _GEN_347 = _T_41 ? _GEN_330 : count; // @[Conditional.scala 39:67 PEArray.scala 101:22]
  wire [2:0] _GEN_348 = _T_41 ? _GEN_331 : state; // @[Conditional.scala 39:67 PEArray.scala 100:22]
  wire [5:0] _GEN_353 = _T_31 ? _GEN_334 : _GEN_346; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_354 = _T_31 ? _GEN_330 : _GEN_347; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_355 = _T_31 ? _GEN_331 : _GEN_348; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_356 = _T_22 ? _GEN_330 : _GEN_354; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_357 = _T_22 ? _GEN_329 : _GEN_353; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_458 = _T_22 ? _GEN_331 : _GEN_355; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_690 = _T_3 ? _GEN_118 : {{2'd0}, GRU_out_width}; // @[Conditional.scala 40:58 PEArray.scala 104:26]
  FP16MulAdder FP16MAC ( // @[PEArray.scala 72:23]
    .io_a(FP16MAC_io_a),
    .io_b(FP16MAC_io_b),
    .io_c(FP16MAC_io_c),
    .io_out(FP16MAC_io_out)
  );
  assign io_ToRightPE = mux3out_reg; // @[PEArray.scala 95:16]
  assign io_ToBelowPE = mux2out_reg; // @[PEArray.scala 94:16]
  assign FP16MAC_io_a = sel1 ? io_FromL1 : io_FromLeftPE; // @[PEArray.scala 50:14 PEArray.scala 50:23 PEArray.scala 51:24]
  assign FP16MAC_io_b = sel5 ? mux4out : _GEN_105; // @[PEArray.scala 77:13 PEArray.scala 78:18 PEArray.scala 81:18]
  assign FP16MAC_io_c = sel5 ? _GEN_105 : mux4out; // @[PEArray.scala 77:13 PEArray.scala 79:18 PEArray.scala 82:18]
  always @(posedge clock) begin
    if (reset) begin // @[PEArray.scala 39:24]
      L0Index <= 6'h0; // @[PEArray.scala 39:24]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h0; // @[PEArray.scala 159:15]
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h9; // @[PEArray.scala 181:15]
      end else begin
        L0Index <= _GEN_357;
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_0 <= _GEN_229;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_1 <= _GEN_230;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_2 <= _GEN_231;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_3 <= _GEN_232;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_4 <= _GEN_233;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_5 <= _GEN_234;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_6 <= _GEN_235;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_7 <= _GEN_236;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_8 <= _GEN_237;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_9 <= _GEN_238;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_10 <= _GEN_239;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_11 <= _GEN_240;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_12 <= _GEN_241;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_13 <= _GEN_242;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_14 <= _GEN_243;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_15 <= _GEN_244;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_16 <= _GEN_245;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_17 <= _GEN_246;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_18 <= _GEN_247;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_19 <= _GEN_248;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_20 <= _GEN_249;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_21 <= _GEN_250;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_22 <= _GEN_251;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_23 <= _GEN_252;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_24 <= _GEN_253;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_25 <= _GEN_254;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_26 <= _GEN_255;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_27 <= _GEN_256;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_28 <= _GEN_257;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_29 <= _GEN_258;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_30 <= _GEN_259;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_31 <= _GEN_260;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_32 <= _GEN_261;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_33 <= _GEN_262;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_34 <= _GEN_263;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_35 <= _GEN_264;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_36 <= _GEN_265;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_37 <= _GEN_266;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_38 <= _GEN_267;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_39 <= _GEN_268;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_40 <= _GEN_269;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_41 <= _GEN_270;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_42 <= _GEN_271;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_43 <= _GEN_272;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_44 <= _GEN_273;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_45 <= _GEN_274;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_46 <= _GEN_275;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_47 <= _GEN_276;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_48 <= _GEN_277;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_49 <= _GEN_278;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_50 <= _GEN_279;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_51 <= _GEN_280;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_52 <= _GEN_281;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_53 <= _GEN_282;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_54 <= _GEN_283;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_55 <= _GEN_284;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_56 <= _GEN_285;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_57 <= _GEN_286;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_58 <= _GEN_287;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_59 <= _GEN_288;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_60 <= _GEN_289;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_61 <= _GEN_290;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_62 <= _GEN_291;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_63 <= _GEN_292;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_64 <= _GEN_293;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_65 <= _GEN_294;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_66 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_67 <= _GEN_296;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_68 <= _GEN_297;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_69 <= _GEN_298;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_70 <= _GEN_299;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_71 <= _GEN_300;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_72 <= _GEN_301;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_73 <= _GEN_302;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_74 <= _GEN_303;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_75 <= _GEN_304;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_76 <= _GEN_305;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_77 <= _GEN_306;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_78 <= _GEN_307;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_79 <= _GEN_308;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_80 <= _GEN_309;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_81 <= _GEN_310;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_82 <= _GEN_311;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_83 <= _GEN_312;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_84 <= _GEN_313;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_85 <= _GEN_314;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_86 <= _GEN_315;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_87 <= _GEN_316;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_88 <= _GEN_317;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_89 <= _GEN_318;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_90 <= _GEN_319;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_91 <= _GEN_320;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_92 <= _GEN_321;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_93 <= _GEN_322;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_94 <= _GEN_323;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_95 <= _GEN_324;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_96 <= _GEN_325;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_97 <= _GEN_326;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_98 <= _GEN_327;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_99 <= _GEN_328;
          end
        end
      end
    end
    if (reset) begin // @[PEArray.scala 100:22]
      state <= 3'h0; // @[PEArray.scala 100:22]
    end else if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[5]) begin // @[PEArray.scala 116:57]
        state <= 3'h1;
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      if (count == 10'h33) begin // @[PEArray.scala 164:27]
        state <= 3'h0; // @[PEArray.scala 166:15]
      end
    end else if (_T_16) begin // @[Conditional.scala 39:67]
      state <= _GEN_126;
    end else begin
      state <= _GEN_458;
    end
    if (reset) begin // @[PEArray.scala 90:28]
      mux2out_reg <= 16'h0; // @[PEArray.scala 90:28]
    end else begin
      mux2out_reg <= MAC_out; // @[PEArray.scala 90:28]
    end
    if (reset) begin // @[PEArray.scala 91:28]
      mux3out_reg <= 16'h0; // @[PEArray.scala 91:28]
    end else if (sel3) begin // @[PEArray.scala 56:14]
      mux3out_reg <= MAC_out; // @[PEArray.scala 56:23]
    end else if (sel1) begin // @[PEArray.scala 50:14]
      mux3out_reg <= io_FromL1; // @[PEArray.scala 50:23]
    end else begin
      mux3out_reg <= io_FromLeftPE; // @[PEArray.scala 51:24]
    end
    if (reset) begin // @[PEArray.scala 101:22]
      count <= 10'h0; // @[PEArray.scala 101:22]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        if (count == 10'h33) begin // @[PEArray.scala 164:27]
          count <= 10'h0; // @[PEArray.scala 165:15]
        end else begin
          count <= _GEN_120;
        end
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        count <= _GEN_125;
      end else begin
        count <= _GEN_356;
      end
    end
    GRU_out_width <= _GEN_690[5:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  L0Index = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  L0Memory_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  L0Memory_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  L0Memory_2 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  L0Memory_3 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  L0Memory_4 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  L0Memory_5 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  L0Memory_6 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  L0Memory_7 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  L0Memory_8 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  L0Memory_9 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  L0Memory_10 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  L0Memory_11 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  L0Memory_12 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  L0Memory_13 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  L0Memory_14 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  L0Memory_15 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  L0Memory_16 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  L0Memory_17 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  L0Memory_18 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  L0Memory_19 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  L0Memory_20 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  L0Memory_21 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  L0Memory_22 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  L0Memory_23 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  L0Memory_24 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  L0Memory_25 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  L0Memory_26 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  L0Memory_27 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  L0Memory_28 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  L0Memory_29 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  L0Memory_30 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  L0Memory_31 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  L0Memory_32 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  L0Memory_33 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  L0Memory_34 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  L0Memory_35 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  L0Memory_36 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  L0Memory_37 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  L0Memory_38 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  L0Memory_39 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  L0Memory_40 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  L0Memory_41 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  L0Memory_42 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  L0Memory_43 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  L0Memory_44 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  L0Memory_45 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  L0Memory_46 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  L0Memory_47 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  L0Memory_48 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  L0Memory_49 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  L0Memory_50 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  L0Memory_51 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  L0Memory_52 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  L0Memory_53 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  L0Memory_54 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  L0Memory_55 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  L0Memory_56 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  L0Memory_57 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  L0Memory_58 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  L0Memory_59 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  L0Memory_60 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  L0Memory_61 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  L0Memory_62 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  L0Memory_63 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  L0Memory_64 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  L0Memory_65 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  L0Memory_66 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  L0Memory_67 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  L0Memory_68 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  L0Memory_69 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  L0Memory_70 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  L0Memory_71 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  L0Memory_72 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  L0Memory_73 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  L0Memory_74 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  L0Memory_75 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  L0Memory_76 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  L0Memory_77 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  L0Memory_78 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  L0Memory_79 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  L0Memory_80 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  L0Memory_81 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  L0Memory_82 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  L0Memory_83 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  L0Memory_84 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  L0Memory_85 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  L0Memory_86 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  L0Memory_87 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  L0Memory_88 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  L0Memory_89 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  L0Memory_90 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  L0Memory_91 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  L0Memory_92 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  L0Memory_93 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  L0Memory_94 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  L0Memory_95 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  L0Memory_96 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  L0Memory_97 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  L0Memory_98 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  L0Memory_99 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  state = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  mux2out_reg = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  mux3out_reg = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  count = _RAND_104[9:0];
  _RAND_105 = {1{`RANDOM}};
  GRU_out_width = _RAND_105[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PE_19(
  input         clock,
  input         reset,
  input  [15:0] io_FromAbovePE,
  input  [15:0] io_FromLeftPE,
  input  [15:0] io_FromL1,
  input  [11:0] io_control_signal_mask,
  output [15:0] io_ToRightPE,
  output [15:0] io_ToBelowPE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] FP16MAC_io_a; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_b; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_c; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_out; // @[PEArray.scala 72:23]
  reg [5:0] L0Index; // @[PEArray.scala 39:24]
  reg [15:0] L0Memory_0; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_1; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_2; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_3; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_4; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_5; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_6; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_7; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_8; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_9; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_10; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_11; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_12; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_13; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_14; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_15; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_16; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_17; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_18; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_19; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_20; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_21; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_22; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_23; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_24; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_25; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_26; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_27; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_28; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_29; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_30; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_31; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_32; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_33; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_34; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_35; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_36; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_37; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_38; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_39; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_40; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_41; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_42; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_43; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_44; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_45; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_46; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_47; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_48; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_49; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_50; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_51; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_52; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_53; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_54; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_55; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_56; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_57; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_58; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_59; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_60; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_61; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_62; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_63; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_64; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_65; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_66; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_67; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_68; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_69; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_70; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_71; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_72; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_73; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_74; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_75; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_76; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_77; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_78; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_79; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_80; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_81; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_82; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_83; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_84; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_85; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_86; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_87; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_88; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_89; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_90; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_91; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_92; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_93; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_94; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_95; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_96; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_97; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_98; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_99; // @[PEArray.scala 40:21]
  reg [2:0] state; // @[PEArray.scala 100:22]
  wire  _T_3 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_12 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_16 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_22 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_31 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_41 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_342 = _T_41 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 231:12 PEArray.scala 32:8]
  wire  _GEN_349 = _T_31 ? 1'h0 : _GEN_342; // @[Conditional.scala 39:67 PEArray.scala 208:12]
  wire  _GEN_459 = _T_22 | _GEN_349; // @[Conditional.scala 39:67 PEArray.scala 32:8]
  wire  _GEN_463 = _T_16 ? 1'h0 : _GEN_459; // @[Conditional.scala 39:67]
  wire  _GEN_572 = _T_12 | _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 149:12]
  wire  sel1 = _T_3 | _GEN_572; // @[Conditional.scala 40:58 PEArray.scala 108:12]
  wire [15:0] MAC_out = FP16MAC_io_out; // @[PEArray.scala 47:21 PEArray.scala 85:11]
  wire  _GEN_465 = _T_16 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 177:12]
  wire  _GEN_580 = _T_12 | _GEN_465; // @[Conditional.scala 39:67 PEArray.scala 34:8]
  wire  sel3 = _T_3 | _GEN_580; // @[Conditional.scala 40:58 PEArray.scala 110:12]
  wire [1:0] _GEN_344 = _T_41 ? 2'h2 : 2'h0; // @[Conditional.scala 39:67 PEArray.scala 233:12 PEArray.scala 35:8]
  wire [1:0] _GEN_351 = _T_31 ? 2'h2 : _GEN_344; // @[Conditional.scala 39:67 PEArray.scala 210:12]
  wire [1:0] _GEN_461 = _T_22 ? 2'h0 : _GEN_351; // @[Conditional.scala 39:67 PEArray.scala 35:8]
  wire [1:0] _GEN_466 = _T_16 ? 2'h0 : _GEN_461; // @[Conditional.scala 39:67 PEArray.scala 178:12]
  wire [1:0] _GEN_574 = _T_12 ? 2'h1 : _GEN_466; // @[Conditional.scala 39:67]
  wire [1:0] sel4 = _T_3 ? 2'h0 : _GEN_574; // @[Conditional.scala 40:58 PEArray.scala 111:12]
  wire [15:0] _GEN_3 = sel4 == 2'h2 ? io_FromL1 : 16'h0; // @[PEArray.scala 65:28 PEArray.scala 66:15 PEArray.scala 69:15]
  wire [15:0] _GEN_4 = sel4 == 2'h1 ? io_FromAbovePE : _GEN_3; // @[PEArray.scala 62:28 PEArray.scala 63:15]
  wire [15:0] mux4out = sel4 == 2'h0 ? 16'h0 : _GEN_4; // @[PEArray.scala 59:22 PEArray.scala 60:13]
  wire [15:0] _GEN_7 = 6'h1 == L0Index ? L0Memory_1 : L0Memory_0; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_8 = 6'h2 == L0Index ? L0Memory_2 : _GEN_7; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_9 = 6'h3 == L0Index ? L0Memory_3 : _GEN_8; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_10 = 6'h4 == L0Index ? L0Memory_4 : _GEN_9; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_11 = 6'h5 == L0Index ? L0Memory_5 : _GEN_10; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_12 = 6'h6 == L0Index ? L0Memory_6 : _GEN_11; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_13 = 6'h7 == L0Index ? L0Memory_7 : _GEN_12; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_14 = 6'h8 == L0Index ? L0Memory_8 : _GEN_13; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_15 = 6'h9 == L0Index ? L0Memory_9 : _GEN_14; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_16 = 6'ha == L0Index ? L0Memory_10 : _GEN_15; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_17 = 6'hb == L0Index ? L0Memory_11 : _GEN_16; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_18 = 6'hc == L0Index ? L0Memory_12 : _GEN_17; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_19 = 6'hd == L0Index ? L0Memory_13 : _GEN_18; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_20 = 6'he == L0Index ? L0Memory_14 : _GEN_19; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_21 = 6'hf == L0Index ? L0Memory_15 : _GEN_20; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_22 = 6'h10 == L0Index ? L0Memory_16 : _GEN_21; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_23 = 6'h11 == L0Index ? L0Memory_17 : _GEN_22; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_24 = 6'h12 == L0Index ? L0Memory_18 : _GEN_23; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_25 = 6'h13 == L0Index ? L0Memory_19 : _GEN_24; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_26 = 6'h14 == L0Index ? L0Memory_20 : _GEN_25; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_27 = 6'h15 == L0Index ? L0Memory_21 : _GEN_26; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_28 = 6'h16 == L0Index ? L0Memory_22 : _GEN_27; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_29 = 6'h17 == L0Index ? L0Memory_23 : _GEN_28; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_30 = 6'h18 == L0Index ? L0Memory_24 : _GEN_29; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_31 = 6'h19 == L0Index ? L0Memory_25 : _GEN_30; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_32 = 6'h1a == L0Index ? L0Memory_26 : _GEN_31; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_33 = 6'h1b == L0Index ? L0Memory_27 : _GEN_32; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_34 = 6'h1c == L0Index ? L0Memory_28 : _GEN_33; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_35 = 6'h1d == L0Index ? L0Memory_29 : _GEN_34; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_36 = 6'h1e == L0Index ? L0Memory_30 : _GEN_35; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_37 = 6'h1f == L0Index ? L0Memory_31 : _GEN_36; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_38 = 6'h20 == L0Index ? L0Memory_32 : _GEN_37; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_39 = 6'h21 == L0Index ? L0Memory_33 : _GEN_38; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_40 = 6'h22 == L0Index ? L0Memory_34 : _GEN_39; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_41 = 6'h23 == L0Index ? L0Memory_35 : _GEN_40; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_42 = 6'h24 == L0Index ? L0Memory_36 : _GEN_41; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_43 = 6'h25 == L0Index ? L0Memory_37 : _GEN_42; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_44 = 6'h26 == L0Index ? L0Memory_38 : _GEN_43; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_45 = 6'h27 == L0Index ? L0Memory_39 : _GEN_44; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_46 = 6'h28 == L0Index ? L0Memory_40 : _GEN_45; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_47 = 6'h29 == L0Index ? L0Memory_41 : _GEN_46; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_48 = 6'h2a == L0Index ? L0Memory_42 : _GEN_47; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_49 = 6'h2b == L0Index ? L0Memory_43 : _GEN_48; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_50 = 6'h2c == L0Index ? L0Memory_44 : _GEN_49; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_51 = 6'h2d == L0Index ? L0Memory_45 : _GEN_50; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_52 = 6'h2e == L0Index ? L0Memory_46 : _GEN_51; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_53 = 6'h2f == L0Index ? L0Memory_47 : _GEN_52; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_54 = 6'h30 == L0Index ? L0Memory_48 : _GEN_53; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_55 = 6'h31 == L0Index ? L0Memory_49 : _GEN_54; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_56 = 6'h32 == L0Index ? L0Memory_50 : _GEN_55; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_57 = 6'h33 == L0Index ? L0Memory_51 : _GEN_56; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_58 = 6'h34 == L0Index ? L0Memory_52 : _GEN_57; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_59 = 6'h35 == L0Index ? L0Memory_53 : _GEN_58; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_60 = 6'h36 == L0Index ? L0Memory_54 : _GEN_59; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_61 = 6'h37 == L0Index ? L0Memory_55 : _GEN_60; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_62 = 6'h38 == L0Index ? L0Memory_56 : _GEN_61; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_63 = 6'h39 == L0Index ? L0Memory_57 : _GEN_62; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_64 = 6'h3a == L0Index ? L0Memory_58 : _GEN_63; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_65 = 6'h3b == L0Index ? L0Memory_59 : _GEN_64; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_66 = 6'h3c == L0Index ? L0Memory_60 : _GEN_65; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_67 = 6'h3d == L0Index ? L0Memory_61 : _GEN_66; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_68 = 6'h3e == L0Index ? L0Memory_62 : _GEN_67; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_69 = 6'h3f == L0Index ? L0Memory_63 : _GEN_68; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [6:0] _GEN_793 = {{1'd0}, L0Index}; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_70 = 7'h40 == _GEN_793 ? L0Memory_64 : _GEN_69; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_71 = 7'h41 == _GEN_793 ? L0Memory_65 : _GEN_70; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_72 = 7'h42 == _GEN_793 ? L0Memory_66 : _GEN_71; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_73 = 7'h43 == _GEN_793 ? L0Memory_67 : _GEN_72; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_74 = 7'h44 == _GEN_793 ? L0Memory_68 : _GEN_73; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_75 = 7'h45 == _GEN_793 ? L0Memory_69 : _GEN_74; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_76 = 7'h46 == _GEN_793 ? L0Memory_70 : _GEN_75; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_77 = 7'h47 == _GEN_793 ? L0Memory_71 : _GEN_76; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_78 = 7'h48 == _GEN_793 ? L0Memory_72 : _GEN_77; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_79 = 7'h49 == _GEN_793 ? L0Memory_73 : _GEN_78; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_80 = 7'h4a == _GEN_793 ? L0Memory_74 : _GEN_79; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_81 = 7'h4b == _GEN_793 ? L0Memory_75 : _GEN_80; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_82 = 7'h4c == _GEN_793 ? L0Memory_76 : _GEN_81; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_83 = 7'h4d == _GEN_793 ? L0Memory_77 : _GEN_82; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_84 = 7'h4e == _GEN_793 ? L0Memory_78 : _GEN_83; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_85 = 7'h4f == _GEN_793 ? L0Memory_79 : _GEN_84; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_86 = 7'h50 == _GEN_793 ? L0Memory_80 : _GEN_85; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_87 = 7'h51 == _GEN_793 ? L0Memory_81 : _GEN_86; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_88 = 7'h52 == _GEN_793 ? L0Memory_82 : _GEN_87; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_89 = 7'h53 == _GEN_793 ? L0Memory_83 : _GEN_88; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_90 = 7'h54 == _GEN_793 ? L0Memory_84 : _GEN_89; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_91 = 7'h55 == _GEN_793 ? L0Memory_85 : _GEN_90; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_92 = 7'h56 == _GEN_793 ? L0Memory_86 : _GEN_91; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_93 = 7'h57 == _GEN_793 ? L0Memory_87 : _GEN_92; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_94 = 7'h58 == _GEN_793 ? L0Memory_88 : _GEN_93; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_95 = 7'h59 == _GEN_793 ? L0Memory_89 : _GEN_94; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_96 = 7'h5a == _GEN_793 ? L0Memory_90 : _GEN_95; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_97 = 7'h5b == _GEN_793 ? L0Memory_91 : _GEN_96; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_98 = 7'h5c == _GEN_793 ? L0Memory_92 : _GEN_97; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_99 = 7'h5d == _GEN_793 ? L0Memory_93 : _GEN_98; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_100 = 7'h5e == _GEN_793 ? L0Memory_94 : _GEN_99; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_101 = 7'h5f == _GEN_793 ? L0Memory_95 : _GEN_100; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_102 = 7'h60 == _GEN_793 ? L0Memory_96 : _GEN_101; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_103 = 7'h61 == _GEN_793 ? L0Memory_97 : _GEN_102; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_104 = 7'h62 == _GEN_793 ? L0Memory_98 : _GEN_103; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_105 = 7'h63 == _GEN_793 ? L0Memory_99 : _GEN_104; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire  _GEN_575 = _T_12 ? 1'h0 : _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 157:12]
  wire  sel5 = _T_3 ? 1'h0 : _GEN_575; // @[Conditional.scala 40:58 PEArray.scala 112:12]
  reg [15:0] mux2out_reg; // @[PEArray.scala 90:28]
  reg [15:0] mux3out_reg; // @[PEArray.scala 91:28]
  reg [9:0] count; // @[PEArray.scala 101:22]
  reg [5:0] GRU_out_width; // @[PEArray.scala 104:26]
  wire [7:0] _GEN_118 = io_control_signal_mask[5] ? 8'h0 : {{2'd0}, GRU_out_width}; // @[PEArray.scala 116:57 PEArray.scala 145:23 PEArray.scala 104:26]
  wire [9:0] _count_T_1 = count + 10'h1; // @[PEArray.scala 162:24]
  wire [9:0] _GEN_120 = count != 10'h33 ? _count_T_1 : count; // @[PEArray.scala 161:27 PEArray.scala 162:15 PEArray.scala 101:22]
  wire [9:0] _GEN_124 = count != 10'h188 ? _count_T_1 : count; // @[PEArray.scala 183:28 PEArray.scala 184:15 PEArray.scala 101:22]
  wire [9:0] _GEN_125 = count == 10'h188 ? 10'h0 : _GEN_124; // @[PEArray.scala 186:28 PEArray.scala 187:15]
  wire [2:0] _GEN_126 = count == 10'h188 ? 3'h0 : state; // @[PEArray.scala 186:28 PEArray.scala 188:15 PEArray.scala 100:22]
  wire [9:0] _GEN_127 = count != 10'h0 ? _count_T_1 : count; // @[PEArray.scala 192:32 PEArray.scala 193:15 PEArray.scala 101:22]
  wire  _T_24 = count == 10'h0; // @[PEArray.scala 195:18]
  wire [5:0] _GEN_128 = count == 10'h0 ? 6'h0 : L0Index; // @[PEArray.scala 195:26 PEArray.scala 196:17 PEArray.scala 39:24]
  wire [9:0] _T_27 = 10'h0 - 10'h1; // @[PEArray.scala 198:51]
  wire [15:0] _GEN_129 = 6'h0 == L0Index ? io_FromL1 : L0Memory_0; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_130 = 6'h1 == L0Index ? io_FromL1 : L0Memory_1; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_131 = 6'h2 == L0Index ? io_FromL1 : L0Memory_2; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_132 = 6'h3 == L0Index ? io_FromL1 : L0Memory_3; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_133 = 6'h4 == L0Index ? io_FromL1 : L0Memory_4; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_134 = 6'h5 == L0Index ? io_FromL1 : L0Memory_5; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_135 = 6'h6 == L0Index ? io_FromL1 : L0Memory_6; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_136 = 6'h7 == L0Index ? io_FromL1 : L0Memory_7; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_137 = 6'h8 == L0Index ? io_FromL1 : L0Memory_8; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_138 = 6'h9 == L0Index ? io_FromL1 : L0Memory_9; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_139 = 6'ha == L0Index ? io_FromL1 : L0Memory_10; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_140 = 6'hb == L0Index ? io_FromL1 : L0Memory_11; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_141 = 6'hc == L0Index ? io_FromL1 : L0Memory_12; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_142 = 6'hd == L0Index ? io_FromL1 : L0Memory_13; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_143 = 6'he == L0Index ? io_FromL1 : L0Memory_14; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_144 = 6'hf == L0Index ? io_FromL1 : L0Memory_15; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_145 = 6'h10 == L0Index ? io_FromL1 : L0Memory_16; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_146 = 6'h11 == L0Index ? io_FromL1 : L0Memory_17; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_147 = 6'h12 == L0Index ? io_FromL1 : L0Memory_18; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_148 = 6'h13 == L0Index ? io_FromL1 : L0Memory_19; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_149 = 6'h14 == L0Index ? io_FromL1 : L0Memory_20; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_150 = 6'h15 == L0Index ? io_FromL1 : L0Memory_21; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_151 = 6'h16 == L0Index ? io_FromL1 : L0Memory_22; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_152 = 6'h17 == L0Index ? io_FromL1 : L0Memory_23; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_153 = 6'h18 == L0Index ? io_FromL1 : L0Memory_24; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_154 = 6'h19 == L0Index ? io_FromL1 : L0Memory_25; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_155 = 6'h1a == L0Index ? io_FromL1 : L0Memory_26; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_156 = 6'h1b == L0Index ? io_FromL1 : L0Memory_27; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_157 = 6'h1c == L0Index ? io_FromL1 : L0Memory_28; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_158 = 6'h1d == L0Index ? io_FromL1 : L0Memory_29; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_159 = 6'h1e == L0Index ? io_FromL1 : L0Memory_30; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_160 = 6'h1f == L0Index ? io_FromL1 : L0Memory_31; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_161 = 6'h20 == L0Index ? io_FromL1 : L0Memory_32; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_162 = 6'h21 == L0Index ? io_FromL1 : L0Memory_33; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_163 = 6'h22 == L0Index ? io_FromL1 : L0Memory_34; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_164 = 6'h23 == L0Index ? io_FromL1 : L0Memory_35; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_165 = 6'h24 == L0Index ? io_FromL1 : L0Memory_36; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_166 = 6'h25 == L0Index ? io_FromL1 : L0Memory_37; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_167 = 6'h26 == L0Index ? io_FromL1 : L0Memory_38; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_168 = 6'h27 == L0Index ? io_FromL1 : L0Memory_39; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_169 = 6'h28 == L0Index ? io_FromL1 : L0Memory_40; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_170 = 6'h29 == L0Index ? io_FromL1 : L0Memory_41; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_171 = 6'h2a == L0Index ? io_FromL1 : L0Memory_42; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_172 = 6'h2b == L0Index ? io_FromL1 : L0Memory_43; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_173 = 6'h2c == L0Index ? io_FromL1 : L0Memory_44; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_174 = 6'h2d == L0Index ? io_FromL1 : L0Memory_45; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_175 = 6'h2e == L0Index ? io_FromL1 : L0Memory_46; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_176 = 6'h2f == L0Index ? io_FromL1 : L0Memory_47; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_177 = 6'h30 == L0Index ? io_FromL1 : L0Memory_48; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_178 = 6'h31 == L0Index ? io_FromL1 : L0Memory_49; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_179 = 6'h32 == L0Index ? io_FromL1 : L0Memory_50; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_180 = 6'h33 == L0Index ? io_FromL1 : L0Memory_51; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_181 = 6'h34 == L0Index ? io_FromL1 : L0Memory_52; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_182 = 6'h35 == L0Index ? io_FromL1 : L0Memory_53; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_183 = 6'h36 == L0Index ? io_FromL1 : L0Memory_54; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_184 = 6'h37 == L0Index ? io_FromL1 : L0Memory_55; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_185 = 6'h38 == L0Index ? io_FromL1 : L0Memory_56; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_186 = 6'h39 == L0Index ? io_FromL1 : L0Memory_57; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_187 = 6'h3a == L0Index ? io_FromL1 : L0Memory_58; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_188 = 6'h3b == L0Index ? io_FromL1 : L0Memory_59; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_189 = 6'h3c == L0Index ? io_FromL1 : L0Memory_60; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_190 = 6'h3d == L0Index ? io_FromL1 : L0Memory_61; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_191 = 6'h3e == L0Index ? io_FromL1 : L0Memory_62; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_192 = 6'h3f == L0Index ? io_FromL1 : L0Memory_63; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_193 = 7'h40 == _GEN_793 ? io_FromL1 : L0Memory_64; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_194 = 7'h41 == _GEN_793 ? io_FromL1 : L0Memory_65; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_195 = 7'h42 == _GEN_793 ? io_FromL1 : L0Memory_66; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_196 = 7'h43 == _GEN_793 ? io_FromL1 : L0Memory_67; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_197 = 7'h44 == _GEN_793 ? io_FromL1 : L0Memory_68; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_198 = 7'h45 == _GEN_793 ? io_FromL1 : L0Memory_69; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_199 = 7'h46 == _GEN_793 ? io_FromL1 : L0Memory_70; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_200 = 7'h47 == _GEN_793 ? io_FromL1 : L0Memory_71; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_201 = 7'h48 == _GEN_793 ? io_FromL1 : L0Memory_72; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_202 = 7'h49 == _GEN_793 ? io_FromL1 : L0Memory_73; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_203 = 7'h4a == _GEN_793 ? io_FromL1 : L0Memory_74; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_204 = 7'h4b == _GEN_793 ? io_FromL1 : L0Memory_75; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_205 = 7'h4c == _GEN_793 ? io_FromL1 : L0Memory_76; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_206 = 7'h4d == _GEN_793 ? io_FromL1 : L0Memory_77; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_207 = 7'h4e == _GEN_793 ? io_FromL1 : L0Memory_78; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_208 = 7'h4f == _GEN_793 ? io_FromL1 : L0Memory_79; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_209 = 7'h50 == _GEN_793 ? io_FromL1 : L0Memory_80; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_210 = 7'h51 == _GEN_793 ? io_FromL1 : L0Memory_81; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_211 = 7'h52 == _GEN_793 ? io_FromL1 : L0Memory_82; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_212 = 7'h53 == _GEN_793 ? io_FromL1 : L0Memory_83; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_213 = 7'h54 == _GEN_793 ? io_FromL1 : L0Memory_84; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_214 = 7'h55 == _GEN_793 ? io_FromL1 : L0Memory_85; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_215 = 7'h56 == _GEN_793 ? io_FromL1 : L0Memory_86; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_216 = 7'h57 == _GEN_793 ? io_FromL1 : L0Memory_87; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_217 = 7'h58 == _GEN_793 ? io_FromL1 : L0Memory_88; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_218 = 7'h59 == _GEN_793 ? io_FromL1 : L0Memory_89; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_219 = 7'h5a == _GEN_793 ? io_FromL1 : L0Memory_90; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_220 = 7'h5b == _GEN_793 ? io_FromL1 : L0Memory_91; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_221 = 7'h5c == _GEN_793 ? io_FromL1 : L0Memory_92; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_222 = 7'h5d == _GEN_793 ? io_FromL1 : L0Memory_93; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_223 = 7'h5e == _GEN_793 ? io_FromL1 : L0Memory_94; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_224 = 7'h5f == _GEN_793 ? io_FromL1 : L0Memory_95; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_225 = 7'h60 == _GEN_793 ? io_FromL1 : L0Memory_96; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_226 = 7'h61 == _GEN_793 ? io_FromL1 : L0Memory_97; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_227 = 7'h62 == _GEN_793 ? io_FromL1 : L0Memory_98; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_228 = 7'h63 == _GEN_793 ? io_FromL1 : L0Memory_99; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [5:0] _L0Index_T_2 = L0Index + 6'h1; // @[PEArray.scala 200:28]
  wire [15:0] _GEN_229 = count >= 10'h1 & count <= _T_27 ? _GEN_129 : L0Memory_0; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_230 = count >= 10'h1 & count <= _T_27 ? _GEN_130 : L0Memory_1; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_231 = count >= 10'h1 & count <= _T_27 ? _GEN_131 : L0Memory_2; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_232 = count >= 10'h1 & count <= _T_27 ? _GEN_132 : L0Memory_3; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_233 = count >= 10'h1 & count <= _T_27 ? _GEN_133 : L0Memory_4; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_234 = count >= 10'h1 & count <= _T_27 ? _GEN_134 : L0Memory_5; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_235 = count >= 10'h1 & count <= _T_27 ? _GEN_135 : L0Memory_6; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_236 = count >= 10'h1 & count <= _T_27 ? _GEN_136 : L0Memory_7; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_237 = count >= 10'h1 & count <= _T_27 ? _GEN_137 : L0Memory_8; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_238 = count >= 10'h1 & count <= _T_27 ? _GEN_138 : L0Memory_9; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_239 = count >= 10'h1 & count <= _T_27 ? _GEN_139 : L0Memory_10; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_240 = count >= 10'h1 & count <= _T_27 ? _GEN_140 : L0Memory_11; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_241 = count >= 10'h1 & count <= _T_27 ? _GEN_141 : L0Memory_12; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_242 = count >= 10'h1 & count <= _T_27 ? _GEN_142 : L0Memory_13; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_243 = count >= 10'h1 & count <= _T_27 ? _GEN_143 : L0Memory_14; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_244 = count >= 10'h1 & count <= _T_27 ? _GEN_144 : L0Memory_15; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_245 = count >= 10'h1 & count <= _T_27 ? _GEN_145 : L0Memory_16; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_246 = count >= 10'h1 & count <= _T_27 ? _GEN_146 : L0Memory_17; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_247 = count >= 10'h1 & count <= _T_27 ? _GEN_147 : L0Memory_18; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_248 = count >= 10'h1 & count <= _T_27 ? _GEN_148 : L0Memory_19; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_249 = count >= 10'h1 & count <= _T_27 ? _GEN_149 : L0Memory_20; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_250 = count >= 10'h1 & count <= _T_27 ? _GEN_150 : L0Memory_21; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_251 = count >= 10'h1 & count <= _T_27 ? _GEN_151 : L0Memory_22; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_252 = count >= 10'h1 & count <= _T_27 ? _GEN_152 : L0Memory_23; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_253 = count >= 10'h1 & count <= _T_27 ? _GEN_153 : L0Memory_24; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_254 = count >= 10'h1 & count <= _T_27 ? _GEN_154 : L0Memory_25; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_255 = count >= 10'h1 & count <= _T_27 ? _GEN_155 : L0Memory_26; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_256 = count >= 10'h1 & count <= _T_27 ? _GEN_156 : L0Memory_27; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_257 = count >= 10'h1 & count <= _T_27 ? _GEN_157 : L0Memory_28; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_258 = count >= 10'h1 & count <= _T_27 ? _GEN_158 : L0Memory_29; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_259 = count >= 10'h1 & count <= _T_27 ? _GEN_159 : L0Memory_30; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_260 = count >= 10'h1 & count <= _T_27 ? _GEN_160 : L0Memory_31; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_261 = count >= 10'h1 & count <= _T_27 ? _GEN_161 : L0Memory_32; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_262 = count >= 10'h1 & count <= _T_27 ? _GEN_162 : L0Memory_33; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_263 = count >= 10'h1 & count <= _T_27 ? _GEN_163 : L0Memory_34; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_264 = count >= 10'h1 & count <= _T_27 ? _GEN_164 : L0Memory_35; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_265 = count >= 10'h1 & count <= _T_27 ? _GEN_165 : L0Memory_36; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_266 = count >= 10'h1 & count <= _T_27 ? _GEN_166 : L0Memory_37; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_267 = count >= 10'h1 & count <= _T_27 ? _GEN_167 : L0Memory_38; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_268 = count >= 10'h1 & count <= _T_27 ? _GEN_168 : L0Memory_39; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_269 = count >= 10'h1 & count <= _T_27 ? _GEN_169 : L0Memory_40; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_270 = count >= 10'h1 & count <= _T_27 ? _GEN_170 : L0Memory_41; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_271 = count >= 10'h1 & count <= _T_27 ? _GEN_171 : L0Memory_42; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_272 = count >= 10'h1 & count <= _T_27 ? _GEN_172 : L0Memory_43; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_273 = count >= 10'h1 & count <= _T_27 ? _GEN_173 : L0Memory_44; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_274 = count >= 10'h1 & count <= _T_27 ? _GEN_174 : L0Memory_45; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_275 = count >= 10'h1 & count <= _T_27 ? _GEN_175 : L0Memory_46; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_276 = count >= 10'h1 & count <= _T_27 ? _GEN_176 : L0Memory_47; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_277 = count >= 10'h1 & count <= _T_27 ? _GEN_177 : L0Memory_48; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_278 = count >= 10'h1 & count <= _T_27 ? _GEN_178 : L0Memory_49; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_279 = count >= 10'h1 & count <= _T_27 ? _GEN_179 : L0Memory_50; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_280 = count >= 10'h1 & count <= _T_27 ? _GEN_180 : L0Memory_51; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_281 = count >= 10'h1 & count <= _T_27 ? _GEN_181 : L0Memory_52; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_282 = count >= 10'h1 & count <= _T_27 ? _GEN_182 : L0Memory_53; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_283 = count >= 10'h1 & count <= _T_27 ? _GEN_183 : L0Memory_54; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_284 = count >= 10'h1 & count <= _T_27 ? _GEN_184 : L0Memory_55; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_285 = count >= 10'h1 & count <= _T_27 ? _GEN_185 : L0Memory_56; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_286 = count >= 10'h1 & count <= _T_27 ? _GEN_186 : L0Memory_57; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_287 = count >= 10'h1 & count <= _T_27 ? _GEN_187 : L0Memory_58; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_288 = count >= 10'h1 & count <= _T_27 ? _GEN_188 : L0Memory_59; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_289 = count >= 10'h1 & count <= _T_27 ? _GEN_189 : L0Memory_60; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_290 = count >= 10'h1 & count <= _T_27 ? _GEN_190 : L0Memory_61; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_291 = count >= 10'h1 & count <= _T_27 ? _GEN_191 : L0Memory_62; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_292 = count >= 10'h1 & count <= _T_27 ? _GEN_192 : L0Memory_63; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_293 = count >= 10'h1 & count <= _T_27 ? _GEN_193 : L0Memory_64; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_294 = count >= 10'h1 & count <= _T_27 ? _GEN_194 : L0Memory_65; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_295 = count >= 10'h1 & count <= _T_27 ? _GEN_195 : L0Memory_66; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_296 = count >= 10'h1 & count <= _T_27 ? _GEN_196 : L0Memory_67; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_297 = count >= 10'h1 & count <= _T_27 ? _GEN_197 : L0Memory_68; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_298 = count >= 10'h1 & count <= _T_27 ? _GEN_198 : L0Memory_69; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_299 = count >= 10'h1 & count <= _T_27 ? _GEN_199 : L0Memory_70; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_300 = count >= 10'h1 & count <= _T_27 ? _GEN_200 : L0Memory_71; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_301 = count >= 10'h1 & count <= _T_27 ? _GEN_201 : L0Memory_72; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_302 = count >= 10'h1 & count <= _T_27 ? _GEN_202 : L0Memory_73; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_303 = count >= 10'h1 & count <= _T_27 ? _GEN_203 : L0Memory_74; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_304 = count >= 10'h1 & count <= _T_27 ? _GEN_204 : L0Memory_75; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_305 = count >= 10'h1 & count <= _T_27 ? _GEN_205 : L0Memory_76; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_306 = count >= 10'h1 & count <= _T_27 ? _GEN_206 : L0Memory_77; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_307 = count >= 10'h1 & count <= _T_27 ? _GEN_207 : L0Memory_78; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_308 = count >= 10'h1 & count <= _T_27 ? _GEN_208 : L0Memory_79; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_309 = count >= 10'h1 & count <= _T_27 ? _GEN_209 : L0Memory_80; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_310 = count >= 10'h1 & count <= _T_27 ? _GEN_210 : L0Memory_81; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_311 = count >= 10'h1 & count <= _T_27 ? _GEN_211 : L0Memory_82; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_312 = count >= 10'h1 & count <= _T_27 ? _GEN_212 : L0Memory_83; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_313 = count >= 10'h1 & count <= _T_27 ? _GEN_213 : L0Memory_84; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_314 = count >= 10'h1 & count <= _T_27 ? _GEN_214 : L0Memory_85; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_315 = count >= 10'h1 & count <= _T_27 ? _GEN_215 : L0Memory_86; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_316 = count >= 10'h1 & count <= _T_27 ? _GEN_216 : L0Memory_87; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_317 = count >= 10'h1 & count <= _T_27 ? _GEN_217 : L0Memory_88; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_318 = count >= 10'h1 & count <= _T_27 ? _GEN_218 : L0Memory_89; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_319 = count >= 10'h1 & count <= _T_27 ? _GEN_219 : L0Memory_90; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_320 = count >= 10'h1 & count <= _T_27 ? _GEN_220 : L0Memory_91; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_321 = count >= 10'h1 & count <= _T_27 ? _GEN_221 : L0Memory_92; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_322 = count >= 10'h1 & count <= _T_27 ? _GEN_222 : L0Memory_93; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_323 = count >= 10'h1 & count <= _T_27 ? _GEN_223 : L0Memory_94; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_324 = count >= 10'h1 & count <= _T_27 ? _GEN_224 : L0Memory_95; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_325 = count >= 10'h1 & count <= _T_27 ? _GEN_225 : L0Memory_96; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_326 = count >= 10'h1 & count <= _T_27 ? _GEN_226 : L0Memory_97; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_327 = count >= 10'h1 & count <= _T_27 ? _GEN_227 : L0Memory_98; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_328 = count >= 10'h1 & count <= _T_27 ? _GEN_228 : L0Memory_99; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [5:0] _GEN_329 = count >= 10'h1 & count <= _T_27 ? _L0Index_T_2 : _GEN_128; // @[PEArray.scala 198:59 PEArray.scala 200:17]
  wire [9:0] _GEN_330 = _T_24 ? 10'h0 : _GEN_127; // @[PEArray.scala 202:32 PEArray.scala 203:15]
  wire [2:0] _GEN_331 = _T_24 ? 3'h0 : state; // @[PEArray.scala 202:32 PEArray.scala 204:15 PEArray.scala 100:22]
  wire [9:0] _GEN_865 = {{4'd0}, GRU_out_width}; // @[PEArray.scala 220:19]
  wire [9:0] _GEN_0 = count % _GEN_865; // @[PEArray.scala 220:19]
  wire [5:0] _T_36 = _GEN_0[5:0]; // @[PEArray.scala 220:19]
  wire [5:0] _T_38 = GRU_out_width - 6'h1; // @[PEArray.scala 220:55]
  wire [5:0] _GEN_334 = _T_36 == _T_38 ? _L0Index_T_2 : 6'h0; // @[PEArray.scala 220:62 PEArray.scala 221:17 PEArray.scala 214:15]
  wire [5:0] _GEN_346 = _T_41 ? _GEN_334 : L0Index; // @[Conditional.scala 39:67 PEArray.scala 39:24]
  wire [9:0] _GEN_347 = _T_41 ? _GEN_330 : count; // @[Conditional.scala 39:67 PEArray.scala 101:22]
  wire [2:0] _GEN_348 = _T_41 ? _GEN_331 : state; // @[Conditional.scala 39:67 PEArray.scala 100:22]
  wire [5:0] _GEN_353 = _T_31 ? _GEN_334 : _GEN_346; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_354 = _T_31 ? _GEN_330 : _GEN_347; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_355 = _T_31 ? _GEN_331 : _GEN_348; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_356 = _T_22 ? _GEN_330 : _GEN_354; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_357 = _T_22 ? _GEN_329 : _GEN_353; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_458 = _T_22 ? _GEN_331 : _GEN_355; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_690 = _T_3 ? _GEN_118 : {{2'd0}, GRU_out_width}; // @[Conditional.scala 40:58 PEArray.scala 104:26]
  FP16MulAdder FP16MAC ( // @[PEArray.scala 72:23]
    .io_a(FP16MAC_io_a),
    .io_b(FP16MAC_io_b),
    .io_c(FP16MAC_io_c),
    .io_out(FP16MAC_io_out)
  );
  assign io_ToRightPE = mux3out_reg; // @[PEArray.scala 95:16]
  assign io_ToBelowPE = mux2out_reg; // @[PEArray.scala 94:16]
  assign FP16MAC_io_a = sel1 ? io_FromL1 : io_FromLeftPE; // @[PEArray.scala 50:14 PEArray.scala 50:23 PEArray.scala 51:24]
  assign FP16MAC_io_b = sel5 ? mux4out : _GEN_105; // @[PEArray.scala 77:13 PEArray.scala 78:18 PEArray.scala 81:18]
  assign FP16MAC_io_c = sel5 ? _GEN_105 : mux4out; // @[PEArray.scala 77:13 PEArray.scala 79:18 PEArray.scala 82:18]
  always @(posedge clock) begin
    if (reset) begin // @[PEArray.scala 39:24]
      L0Index <= 6'h0; // @[PEArray.scala 39:24]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h1; // @[PEArray.scala 159:15]
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h9; // @[PEArray.scala 181:15]
      end else begin
        L0Index <= _GEN_357;
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_0 <= _GEN_229;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_1 <= _GEN_230;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_2 <= _GEN_231;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_3 <= _GEN_232;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_4 <= _GEN_233;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_5 <= _GEN_234;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_6 <= _GEN_235;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_7 <= _GEN_236;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_8 <= _GEN_237;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_9 <= _GEN_238;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_10 <= _GEN_239;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_11 <= _GEN_240;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_12 <= _GEN_241;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_13 <= _GEN_242;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_14 <= _GEN_243;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_15 <= _GEN_244;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_16 <= _GEN_245;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_17 <= _GEN_246;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_18 <= _GEN_247;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_19 <= _GEN_248;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_20 <= _GEN_249;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_21 <= _GEN_250;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_22 <= _GEN_251;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_23 <= _GEN_252;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_24 <= _GEN_253;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_25 <= _GEN_254;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_26 <= _GEN_255;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_27 <= _GEN_256;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_28 <= _GEN_257;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_29 <= _GEN_258;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_30 <= _GEN_259;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_31 <= _GEN_260;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_32 <= _GEN_261;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_33 <= _GEN_262;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_34 <= _GEN_263;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_35 <= _GEN_264;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_36 <= _GEN_265;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_37 <= _GEN_266;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_38 <= _GEN_267;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_39 <= _GEN_268;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_40 <= _GEN_269;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_41 <= _GEN_270;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_42 <= _GEN_271;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_43 <= _GEN_272;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_44 <= _GEN_273;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_45 <= _GEN_274;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_46 <= _GEN_275;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_47 <= _GEN_276;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_48 <= _GEN_277;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_49 <= _GEN_278;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_50 <= _GEN_279;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_51 <= _GEN_280;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_52 <= _GEN_281;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_53 <= _GEN_282;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_54 <= _GEN_283;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_55 <= _GEN_284;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_56 <= _GEN_285;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_57 <= _GEN_286;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_58 <= _GEN_287;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_59 <= _GEN_288;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_60 <= _GEN_289;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_61 <= _GEN_290;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_62 <= _GEN_291;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_63 <= _GEN_292;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_64 <= _GEN_293;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_65 <= _GEN_294;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_66 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_67 <= _GEN_296;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_68 <= _GEN_297;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_69 <= _GEN_298;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_70 <= _GEN_299;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_71 <= _GEN_300;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_72 <= _GEN_301;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_73 <= _GEN_302;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_74 <= _GEN_303;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_75 <= _GEN_304;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_76 <= _GEN_305;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_77 <= _GEN_306;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_78 <= _GEN_307;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_79 <= _GEN_308;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_80 <= _GEN_309;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_81 <= _GEN_310;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_82 <= _GEN_311;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_83 <= _GEN_312;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_84 <= _GEN_313;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_85 <= _GEN_314;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_86 <= _GEN_315;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_87 <= _GEN_316;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_88 <= _GEN_317;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_89 <= _GEN_318;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_90 <= _GEN_319;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_91 <= _GEN_320;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_92 <= _GEN_321;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_93 <= _GEN_322;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_94 <= _GEN_323;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_95 <= _GEN_324;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_96 <= _GEN_325;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_97 <= _GEN_326;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_98 <= _GEN_327;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_99 <= _GEN_328;
          end
        end
      end
    end
    if (reset) begin // @[PEArray.scala 100:22]
      state <= 3'h0; // @[PEArray.scala 100:22]
    end else if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[5]) begin // @[PEArray.scala 116:57]
        state <= 3'h1;
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      if (count == 10'h33) begin // @[PEArray.scala 164:27]
        state <= 3'h0; // @[PEArray.scala 166:15]
      end
    end else if (_T_16) begin // @[Conditional.scala 39:67]
      state <= _GEN_126;
    end else begin
      state <= _GEN_458;
    end
    if (reset) begin // @[PEArray.scala 90:28]
      mux2out_reg <= 16'h0; // @[PEArray.scala 90:28]
    end else begin
      mux2out_reg <= MAC_out; // @[PEArray.scala 90:28]
    end
    if (reset) begin // @[PEArray.scala 91:28]
      mux3out_reg <= 16'h0; // @[PEArray.scala 91:28]
    end else if (sel3) begin // @[PEArray.scala 56:14]
      mux3out_reg <= MAC_out; // @[PEArray.scala 56:23]
    end else if (sel1) begin // @[PEArray.scala 50:14]
      mux3out_reg <= io_FromL1; // @[PEArray.scala 50:23]
    end else begin
      mux3out_reg <= io_FromLeftPE; // @[PEArray.scala 51:24]
    end
    if (reset) begin // @[PEArray.scala 101:22]
      count <= 10'h0; // @[PEArray.scala 101:22]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        if (count == 10'h33) begin // @[PEArray.scala 164:27]
          count <= 10'h0; // @[PEArray.scala 165:15]
        end else begin
          count <= _GEN_120;
        end
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        count <= _GEN_125;
      end else begin
        count <= _GEN_356;
      end
    end
    GRU_out_width <= _GEN_690[5:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  L0Index = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  L0Memory_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  L0Memory_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  L0Memory_2 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  L0Memory_3 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  L0Memory_4 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  L0Memory_5 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  L0Memory_6 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  L0Memory_7 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  L0Memory_8 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  L0Memory_9 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  L0Memory_10 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  L0Memory_11 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  L0Memory_12 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  L0Memory_13 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  L0Memory_14 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  L0Memory_15 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  L0Memory_16 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  L0Memory_17 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  L0Memory_18 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  L0Memory_19 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  L0Memory_20 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  L0Memory_21 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  L0Memory_22 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  L0Memory_23 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  L0Memory_24 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  L0Memory_25 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  L0Memory_26 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  L0Memory_27 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  L0Memory_28 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  L0Memory_29 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  L0Memory_30 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  L0Memory_31 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  L0Memory_32 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  L0Memory_33 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  L0Memory_34 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  L0Memory_35 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  L0Memory_36 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  L0Memory_37 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  L0Memory_38 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  L0Memory_39 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  L0Memory_40 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  L0Memory_41 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  L0Memory_42 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  L0Memory_43 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  L0Memory_44 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  L0Memory_45 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  L0Memory_46 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  L0Memory_47 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  L0Memory_48 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  L0Memory_49 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  L0Memory_50 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  L0Memory_51 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  L0Memory_52 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  L0Memory_53 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  L0Memory_54 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  L0Memory_55 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  L0Memory_56 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  L0Memory_57 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  L0Memory_58 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  L0Memory_59 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  L0Memory_60 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  L0Memory_61 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  L0Memory_62 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  L0Memory_63 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  L0Memory_64 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  L0Memory_65 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  L0Memory_66 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  L0Memory_67 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  L0Memory_68 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  L0Memory_69 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  L0Memory_70 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  L0Memory_71 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  L0Memory_72 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  L0Memory_73 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  L0Memory_74 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  L0Memory_75 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  L0Memory_76 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  L0Memory_77 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  L0Memory_78 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  L0Memory_79 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  L0Memory_80 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  L0Memory_81 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  L0Memory_82 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  L0Memory_83 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  L0Memory_84 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  L0Memory_85 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  L0Memory_86 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  L0Memory_87 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  L0Memory_88 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  L0Memory_89 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  L0Memory_90 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  L0Memory_91 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  L0Memory_92 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  L0Memory_93 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  L0Memory_94 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  L0Memory_95 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  L0Memory_96 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  L0Memory_97 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  L0Memory_98 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  L0Memory_99 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  state = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  mux2out_reg = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  mux3out_reg = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  count = _RAND_104[9:0];
  _RAND_105 = {1{`RANDOM}};
  GRU_out_width = _RAND_105[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PE_20(
  input         clock,
  input         reset,
  input  [15:0] io_FromAbovePE,
  input  [15:0] io_FromLeftPE,
  input  [15:0] io_FromL1,
  input  [2:0]  io_control_signal_control,
  input  [9:0]  io_control_signal_count,
  input  [5:0]  io_control_signal_L0index,
  input  [11:0] io_control_signal_mask,
  input  [7:0]  io_control_signal_gru_out_width,
  output [15:0] io_ToRightPE,
  output [15:0] io_ToBelowPE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] FP16MAC_io_a; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_b; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_c; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_out; // @[PEArray.scala 72:23]
  reg [5:0] L0Index; // @[PEArray.scala 39:24]
  reg [15:0] L0Memory_0; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_1; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_2; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_3; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_4; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_5; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_6; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_7; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_8; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_9; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_10; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_11; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_12; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_13; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_14; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_15; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_16; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_17; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_18; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_19; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_20; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_21; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_22; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_23; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_24; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_25; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_26; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_27; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_28; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_29; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_30; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_31; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_32; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_33; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_34; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_35; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_36; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_37; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_38; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_39; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_40; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_41; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_42; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_43; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_44; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_45; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_46; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_47; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_48; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_49; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_50; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_51; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_52; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_53; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_54; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_55; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_56; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_57; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_58; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_59; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_60; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_61; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_62; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_63; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_64; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_65; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_66; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_67; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_68; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_69; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_70; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_71; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_72; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_73; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_74; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_75; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_76; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_77; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_78; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_79; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_80; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_81; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_82; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_83; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_84; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_85; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_86; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_87; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_88; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_89; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_90; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_91; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_92; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_93; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_94; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_95; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_96; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_97; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_98; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_99; // @[PEArray.scala 40:21]
  reg [2:0] state; // @[PEArray.scala 100:22]
  wire  _T_3 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_12 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_16 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_22 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_31 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_41 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_342 = _T_41 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 231:12 PEArray.scala 32:8]
  wire  _GEN_349 = _T_31 ? 1'h0 : _GEN_342; // @[Conditional.scala 39:67 PEArray.scala 208:12]
  wire  _GEN_459 = _T_22 | _GEN_349; // @[Conditional.scala 39:67 PEArray.scala 32:8]
  wire  _GEN_463 = _T_16 ? 1'h0 : _GEN_459; // @[Conditional.scala 39:67]
  wire  _GEN_572 = _T_12 | _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 149:12]
  wire  sel1 = _T_3 | _GEN_572; // @[Conditional.scala 40:58 PEArray.scala 108:12]
  wire [15:0] MAC_out = FP16MAC_io_out; // @[PEArray.scala 47:21 PEArray.scala 85:11]
  wire  _GEN_465 = _T_16 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 177:12]
  wire  _GEN_580 = _T_12 | _GEN_465; // @[Conditional.scala 39:67 PEArray.scala 34:8]
  wire  sel3 = _T_3 | _GEN_580; // @[Conditional.scala 40:58 PEArray.scala 110:12]
  wire [1:0] _GEN_344 = _T_41 ? 2'h2 : 2'h0; // @[Conditional.scala 39:67 PEArray.scala 233:12 PEArray.scala 35:8]
  wire [1:0] _GEN_351 = _T_31 ? 2'h2 : _GEN_344; // @[Conditional.scala 39:67 PEArray.scala 210:12]
  wire [1:0] _GEN_461 = _T_22 ? 2'h0 : _GEN_351; // @[Conditional.scala 39:67 PEArray.scala 35:8]
  wire [1:0] _GEN_466 = _T_16 ? 2'h0 : _GEN_461; // @[Conditional.scala 39:67 PEArray.scala 178:12]
  wire [1:0] _GEN_574 = _T_12 ? 2'h1 : _GEN_466; // @[Conditional.scala 39:67]
  wire [1:0] sel4 = _T_3 ? 2'h0 : _GEN_574; // @[Conditional.scala 40:58 PEArray.scala 111:12]
  wire [15:0] _GEN_3 = sel4 == 2'h2 ? io_FromL1 : 16'h0; // @[PEArray.scala 65:28 PEArray.scala 66:15 PEArray.scala 69:15]
  wire [15:0] _GEN_4 = sel4 == 2'h1 ? io_FromAbovePE : _GEN_3; // @[PEArray.scala 62:28 PEArray.scala 63:15]
  wire [15:0] mux4out = sel4 == 2'h0 ? 16'h0 : _GEN_4; // @[PEArray.scala 59:22 PEArray.scala 60:13]
  wire [15:0] _GEN_7 = 6'h1 == L0Index ? L0Memory_1 : L0Memory_0; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_8 = 6'h2 == L0Index ? L0Memory_2 : _GEN_7; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_9 = 6'h3 == L0Index ? L0Memory_3 : _GEN_8; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_10 = 6'h4 == L0Index ? L0Memory_4 : _GEN_9; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_11 = 6'h5 == L0Index ? L0Memory_5 : _GEN_10; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_12 = 6'h6 == L0Index ? L0Memory_6 : _GEN_11; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_13 = 6'h7 == L0Index ? L0Memory_7 : _GEN_12; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_14 = 6'h8 == L0Index ? L0Memory_8 : _GEN_13; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_15 = 6'h9 == L0Index ? L0Memory_9 : _GEN_14; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_16 = 6'ha == L0Index ? L0Memory_10 : _GEN_15; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_17 = 6'hb == L0Index ? L0Memory_11 : _GEN_16; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_18 = 6'hc == L0Index ? L0Memory_12 : _GEN_17; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_19 = 6'hd == L0Index ? L0Memory_13 : _GEN_18; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_20 = 6'he == L0Index ? L0Memory_14 : _GEN_19; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_21 = 6'hf == L0Index ? L0Memory_15 : _GEN_20; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_22 = 6'h10 == L0Index ? L0Memory_16 : _GEN_21; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_23 = 6'h11 == L0Index ? L0Memory_17 : _GEN_22; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_24 = 6'h12 == L0Index ? L0Memory_18 : _GEN_23; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_25 = 6'h13 == L0Index ? L0Memory_19 : _GEN_24; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_26 = 6'h14 == L0Index ? L0Memory_20 : _GEN_25; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_27 = 6'h15 == L0Index ? L0Memory_21 : _GEN_26; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_28 = 6'h16 == L0Index ? L0Memory_22 : _GEN_27; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_29 = 6'h17 == L0Index ? L0Memory_23 : _GEN_28; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_30 = 6'h18 == L0Index ? L0Memory_24 : _GEN_29; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_31 = 6'h19 == L0Index ? L0Memory_25 : _GEN_30; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_32 = 6'h1a == L0Index ? L0Memory_26 : _GEN_31; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_33 = 6'h1b == L0Index ? L0Memory_27 : _GEN_32; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_34 = 6'h1c == L0Index ? L0Memory_28 : _GEN_33; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_35 = 6'h1d == L0Index ? L0Memory_29 : _GEN_34; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_36 = 6'h1e == L0Index ? L0Memory_30 : _GEN_35; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_37 = 6'h1f == L0Index ? L0Memory_31 : _GEN_36; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_38 = 6'h20 == L0Index ? L0Memory_32 : _GEN_37; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_39 = 6'h21 == L0Index ? L0Memory_33 : _GEN_38; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_40 = 6'h22 == L0Index ? L0Memory_34 : _GEN_39; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_41 = 6'h23 == L0Index ? L0Memory_35 : _GEN_40; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_42 = 6'h24 == L0Index ? L0Memory_36 : _GEN_41; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_43 = 6'h25 == L0Index ? L0Memory_37 : _GEN_42; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_44 = 6'h26 == L0Index ? L0Memory_38 : _GEN_43; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_45 = 6'h27 == L0Index ? L0Memory_39 : _GEN_44; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_46 = 6'h28 == L0Index ? L0Memory_40 : _GEN_45; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_47 = 6'h29 == L0Index ? L0Memory_41 : _GEN_46; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_48 = 6'h2a == L0Index ? L0Memory_42 : _GEN_47; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_49 = 6'h2b == L0Index ? L0Memory_43 : _GEN_48; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_50 = 6'h2c == L0Index ? L0Memory_44 : _GEN_49; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_51 = 6'h2d == L0Index ? L0Memory_45 : _GEN_50; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_52 = 6'h2e == L0Index ? L0Memory_46 : _GEN_51; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_53 = 6'h2f == L0Index ? L0Memory_47 : _GEN_52; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_54 = 6'h30 == L0Index ? L0Memory_48 : _GEN_53; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_55 = 6'h31 == L0Index ? L0Memory_49 : _GEN_54; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_56 = 6'h32 == L0Index ? L0Memory_50 : _GEN_55; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_57 = 6'h33 == L0Index ? L0Memory_51 : _GEN_56; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_58 = 6'h34 == L0Index ? L0Memory_52 : _GEN_57; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_59 = 6'h35 == L0Index ? L0Memory_53 : _GEN_58; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_60 = 6'h36 == L0Index ? L0Memory_54 : _GEN_59; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_61 = 6'h37 == L0Index ? L0Memory_55 : _GEN_60; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_62 = 6'h38 == L0Index ? L0Memory_56 : _GEN_61; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_63 = 6'h39 == L0Index ? L0Memory_57 : _GEN_62; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_64 = 6'h3a == L0Index ? L0Memory_58 : _GEN_63; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_65 = 6'h3b == L0Index ? L0Memory_59 : _GEN_64; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_66 = 6'h3c == L0Index ? L0Memory_60 : _GEN_65; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_67 = 6'h3d == L0Index ? L0Memory_61 : _GEN_66; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_68 = 6'h3e == L0Index ? L0Memory_62 : _GEN_67; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_69 = 6'h3f == L0Index ? L0Memory_63 : _GEN_68; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [6:0] _GEN_793 = {{1'd0}, L0Index}; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_70 = 7'h40 == _GEN_793 ? L0Memory_64 : _GEN_69; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_71 = 7'h41 == _GEN_793 ? L0Memory_65 : _GEN_70; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_72 = 7'h42 == _GEN_793 ? L0Memory_66 : _GEN_71; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_73 = 7'h43 == _GEN_793 ? L0Memory_67 : _GEN_72; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_74 = 7'h44 == _GEN_793 ? L0Memory_68 : _GEN_73; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_75 = 7'h45 == _GEN_793 ? L0Memory_69 : _GEN_74; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_76 = 7'h46 == _GEN_793 ? L0Memory_70 : _GEN_75; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_77 = 7'h47 == _GEN_793 ? L0Memory_71 : _GEN_76; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_78 = 7'h48 == _GEN_793 ? L0Memory_72 : _GEN_77; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_79 = 7'h49 == _GEN_793 ? L0Memory_73 : _GEN_78; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_80 = 7'h4a == _GEN_793 ? L0Memory_74 : _GEN_79; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_81 = 7'h4b == _GEN_793 ? L0Memory_75 : _GEN_80; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_82 = 7'h4c == _GEN_793 ? L0Memory_76 : _GEN_81; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_83 = 7'h4d == _GEN_793 ? L0Memory_77 : _GEN_82; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_84 = 7'h4e == _GEN_793 ? L0Memory_78 : _GEN_83; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_85 = 7'h4f == _GEN_793 ? L0Memory_79 : _GEN_84; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_86 = 7'h50 == _GEN_793 ? L0Memory_80 : _GEN_85; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_87 = 7'h51 == _GEN_793 ? L0Memory_81 : _GEN_86; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_88 = 7'h52 == _GEN_793 ? L0Memory_82 : _GEN_87; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_89 = 7'h53 == _GEN_793 ? L0Memory_83 : _GEN_88; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_90 = 7'h54 == _GEN_793 ? L0Memory_84 : _GEN_89; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_91 = 7'h55 == _GEN_793 ? L0Memory_85 : _GEN_90; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_92 = 7'h56 == _GEN_793 ? L0Memory_86 : _GEN_91; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_93 = 7'h57 == _GEN_793 ? L0Memory_87 : _GEN_92; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_94 = 7'h58 == _GEN_793 ? L0Memory_88 : _GEN_93; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_95 = 7'h59 == _GEN_793 ? L0Memory_89 : _GEN_94; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_96 = 7'h5a == _GEN_793 ? L0Memory_90 : _GEN_95; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_97 = 7'h5b == _GEN_793 ? L0Memory_91 : _GEN_96; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_98 = 7'h5c == _GEN_793 ? L0Memory_92 : _GEN_97; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_99 = 7'h5d == _GEN_793 ? L0Memory_93 : _GEN_98; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_100 = 7'h5e == _GEN_793 ? L0Memory_94 : _GEN_99; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_101 = 7'h5f == _GEN_793 ? L0Memory_95 : _GEN_100; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_102 = 7'h60 == _GEN_793 ? L0Memory_96 : _GEN_101; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_103 = 7'h61 == _GEN_793 ? L0Memory_97 : _GEN_102; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_104 = 7'h62 == _GEN_793 ? L0Memory_98 : _GEN_103; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_105 = 7'h63 == _GEN_793 ? L0Memory_99 : _GEN_104; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire  _GEN_575 = _T_12 ? 1'h0 : _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 157:12]
  wire  sel5 = _T_3 ? 1'h0 : _GEN_575; // @[Conditional.scala 40:58 PEArray.scala 112:12]
  reg [15:0] mux2out_reg; // @[PEArray.scala 90:28]
  reg [15:0] mux3out_reg; // @[PEArray.scala 91:28]
  reg [9:0] count; // @[PEArray.scala 101:22]
  reg [9:0] count_max; // @[PEArray.scala 102:22]
  reg [5:0] L0index_begin; // @[PEArray.scala 103:26]
  reg [5:0] GRU_out_width; // @[PEArray.scala 104:26]
  wire  _T_6 = 3'h0 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_7 = 3'h1 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_8 = 3'h2 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_9 = 3'h3 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_10 = 3'h4 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_11 = 3'h5 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_109 = _T_11 ? 3'h5 : state; // @[Conditional.scala 39:67 PEArray.scala 140:19 PEArray.scala 100:22]
  wire [2:0] _GEN_110 = _T_10 ? 3'h4 : _GEN_109; // @[Conditional.scala 39:67 PEArray.scala 136:19]
  wire [2:0] _GEN_111 = _T_9 ? 3'h3 : _GEN_110; // @[Conditional.scala 39:67 PEArray.scala 132:19]
  wire [2:0] _GEN_112 = _T_8 ? 3'h2 : _GEN_111; // @[Conditional.scala 39:67 PEArray.scala 128:19]
  wire [2:0] _GEN_113 = _T_7 ? 3'h1 : _GEN_112; // @[Conditional.scala 39:67 PEArray.scala 124:19]
  wire [7:0] _GEN_118 = io_control_signal_mask[5] ? io_control_signal_gru_out_width : {{2'd0}, GRU_out_width}; // @[PEArray.scala 116:57 PEArray.scala 145:23 PEArray.scala 104:26]
  wire [9:0] _count_T_1 = count + 10'h1; // @[PEArray.scala 162:24]
  wire [9:0] _GEN_120 = count != 10'h33 ? _count_T_1 : count; // @[PEArray.scala 161:27 PEArray.scala 162:15 PEArray.scala 101:22]
  wire [9:0] _GEN_124 = count != 10'h188 ? _count_T_1 : count; // @[PEArray.scala 183:28 PEArray.scala 184:15 PEArray.scala 101:22]
  wire [9:0] _GEN_125 = count == 10'h188 ? 10'h0 : _GEN_124; // @[PEArray.scala 186:28 PEArray.scala 187:15]
  wire [2:0] _GEN_126 = count == 10'h188 ? 3'h0 : state; // @[PEArray.scala 186:28 PEArray.scala 188:15 PEArray.scala 100:22]
  wire [9:0] _GEN_127 = count != count_max ? _count_T_1 : count; // @[PEArray.scala 192:32 PEArray.scala 193:15 PEArray.scala 101:22]
  wire [5:0] _GEN_128 = count == 10'h0 ? L0index_begin : L0Index; // @[PEArray.scala 195:26 PEArray.scala 196:17 PEArray.scala 39:24]
  wire [9:0] _T_27 = count_max - 10'h1; // @[PEArray.scala 198:51]
  wire [15:0] _GEN_129 = 6'h0 == L0Index ? io_FromL1 : L0Memory_0; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_130 = 6'h1 == L0Index ? io_FromL1 : L0Memory_1; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_131 = 6'h2 == L0Index ? io_FromL1 : L0Memory_2; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_132 = 6'h3 == L0Index ? io_FromL1 : L0Memory_3; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_133 = 6'h4 == L0Index ? io_FromL1 : L0Memory_4; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_134 = 6'h5 == L0Index ? io_FromL1 : L0Memory_5; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_135 = 6'h6 == L0Index ? io_FromL1 : L0Memory_6; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_136 = 6'h7 == L0Index ? io_FromL1 : L0Memory_7; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_137 = 6'h8 == L0Index ? io_FromL1 : L0Memory_8; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_138 = 6'h9 == L0Index ? io_FromL1 : L0Memory_9; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_139 = 6'ha == L0Index ? io_FromL1 : L0Memory_10; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_140 = 6'hb == L0Index ? io_FromL1 : L0Memory_11; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_141 = 6'hc == L0Index ? io_FromL1 : L0Memory_12; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_142 = 6'hd == L0Index ? io_FromL1 : L0Memory_13; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_143 = 6'he == L0Index ? io_FromL1 : L0Memory_14; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_144 = 6'hf == L0Index ? io_FromL1 : L0Memory_15; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_145 = 6'h10 == L0Index ? io_FromL1 : L0Memory_16; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_146 = 6'h11 == L0Index ? io_FromL1 : L0Memory_17; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_147 = 6'h12 == L0Index ? io_FromL1 : L0Memory_18; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_148 = 6'h13 == L0Index ? io_FromL1 : L0Memory_19; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_149 = 6'h14 == L0Index ? io_FromL1 : L0Memory_20; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_150 = 6'h15 == L0Index ? io_FromL1 : L0Memory_21; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_151 = 6'h16 == L0Index ? io_FromL1 : L0Memory_22; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_152 = 6'h17 == L0Index ? io_FromL1 : L0Memory_23; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_153 = 6'h18 == L0Index ? io_FromL1 : L0Memory_24; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_154 = 6'h19 == L0Index ? io_FromL1 : L0Memory_25; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_155 = 6'h1a == L0Index ? io_FromL1 : L0Memory_26; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_156 = 6'h1b == L0Index ? io_FromL1 : L0Memory_27; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_157 = 6'h1c == L0Index ? io_FromL1 : L0Memory_28; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_158 = 6'h1d == L0Index ? io_FromL1 : L0Memory_29; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_159 = 6'h1e == L0Index ? io_FromL1 : L0Memory_30; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_160 = 6'h1f == L0Index ? io_FromL1 : L0Memory_31; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_161 = 6'h20 == L0Index ? io_FromL1 : L0Memory_32; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_162 = 6'h21 == L0Index ? io_FromL1 : L0Memory_33; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_163 = 6'h22 == L0Index ? io_FromL1 : L0Memory_34; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_164 = 6'h23 == L0Index ? io_FromL1 : L0Memory_35; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_165 = 6'h24 == L0Index ? io_FromL1 : L0Memory_36; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_166 = 6'h25 == L0Index ? io_FromL1 : L0Memory_37; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_167 = 6'h26 == L0Index ? io_FromL1 : L0Memory_38; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_168 = 6'h27 == L0Index ? io_FromL1 : L0Memory_39; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_169 = 6'h28 == L0Index ? io_FromL1 : L0Memory_40; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_170 = 6'h29 == L0Index ? io_FromL1 : L0Memory_41; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_171 = 6'h2a == L0Index ? io_FromL1 : L0Memory_42; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_172 = 6'h2b == L0Index ? io_FromL1 : L0Memory_43; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_173 = 6'h2c == L0Index ? io_FromL1 : L0Memory_44; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_174 = 6'h2d == L0Index ? io_FromL1 : L0Memory_45; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_175 = 6'h2e == L0Index ? io_FromL1 : L0Memory_46; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_176 = 6'h2f == L0Index ? io_FromL1 : L0Memory_47; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_177 = 6'h30 == L0Index ? io_FromL1 : L0Memory_48; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_178 = 6'h31 == L0Index ? io_FromL1 : L0Memory_49; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_179 = 6'h32 == L0Index ? io_FromL1 : L0Memory_50; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_180 = 6'h33 == L0Index ? io_FromL1 : L0Memory_51; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_181 = 6'h34 == L0Index ? io_FromL1 : L0Memory_52; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_182 = 6'h35 == L0Index ? io_FromL1 : L0Memory_53; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_183 = 6'h36 == L0Index ? io_FromL1 : L0Memory_54; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_184 = 6'h37 == L0Index ? io_FromL1 : L0Memory_55; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_185 = 6'h38 == L0Index ? io_FromL1 : L0Memory_56; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_186 = 6'h39 == L0Index ? io_FromL1 : L0Memory_57; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_187 = 6'h3a == L0Index ? io_FromL1 : L0Memory_58; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_188 = 6'h3b == L0Index ? io_FromL1 : L0Memory_59; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_189 = 6'h3c == L0Index ? io_FromL1 : L0Memory_60; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_190 = 6'h3d == L0Index ? io_FromL1 : L0Memory_61; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_191 = 6'h3e == L0Index ? io_FromL1 : L0Memory_62; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_192 = 6'h3f == L0Index ? io_FromL1 : L0Memory_63; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_193 = 7'h40 == _GEN_793 ? io_FromL1 : L0Memory_64; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_194 = 7'h41 == _GEN_793 ? io_FromL1 : L0Memory_65; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_195 = 7'h42 == _GEN_793 ? io_FromL1 : L0Memory_66; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_196 = 7'h43 == _GEN_793 ? io_FromL1 : L0Memory_67; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_197 = 7'h44 == _GEN_793 ? io_FromL1 : L0Memory_68; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_198 = 7'h45 == _GEN_793 ? io_FromL1 : L0Memory_69; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_199 = 7'h46 == _GEN_793 ? io_FromL1 : L0Memory_70; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_200 = 7'h47 == _GEN_793 ? io_FromL1 : L0Memory_71; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_201 = 7'h48 == _GEN_793 ? io_FromL1 : L0Memory_72; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_202 = 7'h49 == _GEN_793 ? io_FromL1 : L0Memory_73; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_203 = 7'h4a == _GEN_793 ? io_FromL1 : L0Memory_74; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_204 = 7'h4b == _GEN_793 ? io_FromL1 : L0Memory_75; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_205 = 7'h4c == _GEN_793 ? io_FromL1 : L0Memory_76; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_206 = 7'h4d == _GEN_793 ? io_FromL1 : L0Memory_77; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_207 = 7'h4e == _GEN_793 ? io_FromL1 : L0Memory_78; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_208 = 7'h4f == _GEN_793 ? io_FromL1 : L0Memory_79; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_209 = 7'h50 == _GEN_793 ? io_FromL1 : L0Memory_80; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_210 = 7'h51 == _GEN_793 ? io_FromL1 : L0Memory_81; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_211 = 7'h52 == _GEN_793 ? io_FromL1 : L0Memory_82; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_212 = 7'h53 == _GEN_793 ? io_FromL1 : L0Memory_83; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_213 = 7'h54 == _GEN_793 ? io_FromL1 : L0Memory_84; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_214 = 7'h55 == _GEN_793 ? io_FromL1 : L0Memory_85; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_215 = 7'h56 == _GEN_793 ? io_FromL1 : L0Memory_86; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_216 = 7'h57 == _GEN_793 ? io_FromL1 : L0Memory_87; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_217 = 7'h58 == _GEN_793 ? io_FromL1 : L0Memory_88; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_218 = 7'h59 == _GEN_793 ? io_FromL1 : L0Memory_89; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_219 = 7'h5a == _GEN_793 ? io_FromL1 : L0Memory_90; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_220 = 7'h5b == _GEN_793 ? io_FromL1 : L0Memory_91; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_221 = 7'h5c == _GEN_793 ? io_FromL1 : L0Memory_92; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_222 = 7'h5d == _GEN_793 ? io_FromL1 : L0Memory_93; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_223 = 7'h5e == _GEN_793 ? io_FromL1 : L0Memory_94; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_224 = 7'h5f == _GEN_793 ? io_FromL1 : L0Memory_95; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_225 = 7'h60 == _GEN_793 ? io_FromL1 : L0Memory_96; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_226 = 7'h61 == _GEN_793 ? io_FromL1 : L0Memory_97; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_227 = 7'h62 == _GEN_793 ? io_FromL1 : L0Memory_98; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_228 = 7'h63 == _GEN_793 ? io_FromL1 : L0Memory_99; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [5:0] _L0Index_T_2 = L0Index + 6'h1; // @[PEArray.scala 200:28]
  wire [15:0] _GEN_229 = count >= 10'h1 & count <= _T_27 ? _GEN_129 : L0Memory_0; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_230 = count >= 10'h1 & count <= _T_27 ? _GEN_130 : L0Memory_1; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_231 = count >= 10'h1 & count <= _T_27 ? _GEN_131 : L0Memory_2; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_232 = count >= 10'h1 & count <= _T_27 ? _GEN_132 : L0Memory_3; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_233 = count >= 10'h1 & count <= _T_27 ? _GEN_133 : L0Memory_4; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_234 = count >= 10'h1 & count <= _T_27 ? _GEN_134 : L0Memory_5; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_235 = count >= 10'h1 & count <= _T_27 ? _GEN_135 : L0Memory_6; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_236 = count >= 10'h1 & count <= _T_27 ? _GEN_136 : L0Memory_7; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_237 = count >= 10'h1 & count <= _T_27 ? _GEN_137 : L0Memory_8; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_238 = count >= 10'h1 & count <= _T_27 ? _GEN_138 : L0Memory_9; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_239 = count >= 10'h1 & count <= _T_27 ? _GEN_139 : L0Memory_10; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_240 = count >= 10'h1 & count <= _T_27 ? _GEN_140 : L0Memory_11; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_241 = count >= 10'h1 & count <= _T_27 ? _GEN_141 : L0Memory_12; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_242 = count >= 10'h1 & count <= _T_27 ? _GEN_142 : L0Memory_13; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_243 = count >= 10'h1 & count <= _T_27 ? _GEN_143 : L0Memory_14; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_244 = count >= 10'h1 & count <= _T_27 ? _GEN_144 : L0Memory_15; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_245 = count >= 10'h1 & count <= _T_27 ? _GEN_145 : L0Memory_16; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_246 = count >= 10'h1 & count <= _T_27 ? _GEN_146 : L0Memory_17; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_247 = count >= 10'h1 & count <= _T_27 ? _GEN_147 : L0Memory_18; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_248 = count >= 10'h1 & count <= _T_27 ? _GEN_148 : L0Memory_19; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_249 = count >= 10'h1 & count <= _T_27 ? _GEN_149 : L0Memory_20; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_250 = count >= 10'h1 & count <= _T_27 ? _GEN_150 : L0Memory_21; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_251 = count >= 10'h1 & count <= _T_27 ? _GEN_151 : L0Memory_22; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_252 = count >= 10'h1 & count <= _T_27 ? _GEN_152 : L0Memory_23; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_253 = count >= 10'h1 & count <= _T_27 ? _GEN_153 : L0Memory_24; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_254 = count >= 10'h1 & count <= _T_27 ? _GEN_154 : L0Memory_25; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_255 = count >= 10'h1 & count <= _T_27 ? _GEN_155 : L0Memory_26; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_256 = count >= 10'h1 & count <= _T_27 ? _GEN_156 : L0Memory_27; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_257 = count >= 10'h1 & count <= _T_27 ? _GEN_157 : L0Memory_28; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_258 = count >= 10'h1 & count <= _T_27 ? _GEN_158 : L0Memory_29; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_259 = count >= 10'h1 & count <= _T_27 ? _GEN_159 : L0Memory_30; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_260 = count >= 10'h1 & count <= _T_27 ? _GEN_160 : L0Memory_31; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_261 = count >= 10'h1 & count <= _T_27 ? _GEN_161 : L0Memory_32; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_262 = count >= 10'h1 & count <= _T_27 ? _GEN_162 : L0Memory_33; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_263 = count >= 10'h1 & count <= _T_27 ? _GEN_163 : L0Memory_34; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_264 = count >= 10'h1 & count <= _T_27 ? _GEN_164 : L0Memory_35; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_265 = count >= 10'h1 & count <= _T_27 ? _GEN_165 : L0Memory_36; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_266 = count >= 10'h1 & count <= _T_27 ? _GEN_166 : L0Memory_37; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_267 = count >= 10'h1 & count <= _T_27 ? _GEN_167 : L0Memory_38; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_268 = count >= 10'h1 & count <= _T_27 ? _GEN_168 : L0Memory_39; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_269 = count >= 10'h1 & count <= _T_27 ? _GEN_169 : L0Memory_40; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_270 = count >= 10'h1 & count <= _T_27 ? _GEN_170 : L0Memory_41; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_271 = count >= 10'h1 & count <= _T_27 ? _GEN_171 : L0Memory_42; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_272 = count >= 10'h1 & count <= _T_27 ? _GEN_172 : L0Memory_43; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_273 = count >= 10'h1 & count <= _T_27 ? _GEN_173 : L0Memory_44; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_274 = count >= 10'h1 & count <= _T_27 ? _GEN_174 : L0Memory_45; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_275 = count >= 10'h1 & count <= _T_27 ? _GEN_175 : L0Memory_46; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_276 = count >= 10'h1 & count <= _T_27 ? _GEN_176 : L0Memory_47; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_277 = count >= 10'h1 & count <= _T_27 ? _GEN_177 : L0Memory_48; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_278 = count >= 10'h1 & count <= _T_27 ? _GEN_178 : L0Memory_49; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_279 = count >= 10'h1 & count <= _T_27 ? _GEN_179 : L0Memory_50; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_280 = count >= 10'h1 & count <= _T_27 ? _GEN_180 : L0Memory_51; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_281 = count >= 10'h1 & count <= _T_27 ? _GEN_181 : L0Memory_52; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_282 = count >= 10'h1 & count <= _T_27 ? _GEN_182 : L0Memory_53; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_283 = count >= 10'h1 & count <= _T_27 ? _GEN_183 : L0Memory_54; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_284 = count >= 10'h1 & count <= _T_27 ? _GEN_184 : L0Memory_55; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_285 = count >= 10'h1 & count <= _T_27 ? _GEN_185 : L0Memory_56; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_286 = count >= 10'h1 & count <= _T_27 ? _GEN_186 : L0Memory_57; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_287 = count >= 10'h1 & count <= _T_27 ? _GEN_187 : L0Memory_58; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_288 = count >= 10'h1 & count <= _T_27 ? _GEN_188 : L0Memory_59; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_289 = count >= 10'h1 & count <= _T_27 ? _GEN_189 : L0Memory_60; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_290 = count >= 10'h1 & count <= _T_27 ? _GEN_190 : L0Memory_61; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_291 = count >= 10'h1 & count <= _T_27 ? _GEN_191 : L0Memory_62; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_292 = count >= 10'h1 & count <= _T_27 ? _GEN_192 : L0Memory_63; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_293 = count >= 10'h1 & count <= _T_27 ? _GEN_193 : L0Memory_64; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_294 = count >= 10'h1 & count <= _T_27 ? _GEN_194 : L0Memory_65; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_295 = count >= 10'h1 & count <= _T_27 ? _GEN_195 : L0Memory_66; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_296 = count >= 10'h1 & count <= _T_27 ? _GEN_196 : L0Memory_67; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_297 = count >= 10'h1 & count <= _T_27 ? _GEN_197 : L0Memory_68; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_298 = count >= 10'h1 & count <= _T_27 ? _GEN_198 : L0Memory_69; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_299 = count >= 10'h1 & count <= _T_27 ? _GEN_199 : L0Memory_70; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_300 = count >= 10'h1 & count <= _T_27 ? _GEN_200 : L0Memory_71; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_301 = count >= 10'h1 & count <= _T_27 ? _GEN_201 : L0Memory_72; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_302 = count >= 10'h1 & count <= _T_27 ? _GEN_202 : L0Memory_73; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_303 = count >= 10'h1 & count <= _T_27 ? _GEN_203 : L0Memory_74; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_304 = count >= 10'h1 & count <= _T_27 ? _GEN_204 : L0Memory_75; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_305 = count >= 10'h1 & count <= _T_27 ? _GEN_205 : L0Memory_76; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_306 = count >= 10'h1 & count <= _T_27 ? _GEN_206 : L0Memory_77; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_307 = count >= 10'h1 & count <= _T_27 ? _GEN_207 : L0Memory_78; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_308 = count >= 10'h1 & count <= _T_27 ? _GEN_208 : L0Memory_79; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_309 = count >= 10'h1 & count <= _T_27 ? _GEN_209 : L0Memory_80; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_310 = count >= 10'h1 & count <= _T_27 ? _GEN_210 : L0Memory_81; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_311 = count >= 10'h1 & count <= _T_27 ? _GEN_211 : L0Memory_82; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_312 = count >= 10'h1 & count <= _T_27 ? _GEN_212 : L0Memory_83; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_313 = count >= 10'h1 & count <= _T_27 ? _GEN_213 : L0Memory_84; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_314 = count >= 10'h1 & count <= _T_27 ? _GEN_214 : L0Memory_85; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_315 = count >= 10'h1 & count <= _T_27 ? _GEN_215 : L0Memory_86; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_316 = count >= 10'h1 & count <= _T_27 ? _GEN_216 : L0Memory_87; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_317 = count >= 10'h1 & count <= _T_27 ? _GEN_217 : L0Memory_88; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_318 = count >= 10'h1 & count <= _T_27 ? _GEN_218 : L0Memory_89; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_319 = count >= 10'h1 & count <= _T_27 ? _GEN_219 : L0Memory_90; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_320 = count >= 10'h1 & count <= _T_27 ? _GEN_220 : L0Memory_91; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_321 = count >= 10'h1 & count <= _T_27 ? _GEN_221 : L0Memory_92; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_322 = count >= 10'h1 & count <= _T_27 ? _GEN_222 : L0Memory_93; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_323 = count >= 10'h1 & count <= _T_27 ? _GEN_223 : L0Memory_94; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_324 = count >= 10'h1 & count <= _T_27 ? _GEN_224 : L0Memory_95; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_325 = count >= 10'h1 & count <= _T_27 ? _GEN_225 : L0Memory_96; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_326 = count >= 10'h1 & count <= _T_27 ? _GEN_226 : L0Memory_97; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_327 = count >= 10'h1 & count <= _T_27 ? _GEN_227 : L0Memory_98; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_328 = count >= 10'h1 & count <= _T_27 ? _GEN_228 : L0Memory_99; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [5:0] _GEN_329 = count >= 10'h1 & count <= _T_27 ? _L0Index_T_2 : _GEN_128; // @[PEArray.scala 198:59 PEArray.scala 200:17]
  wire [9:0] _GEN_330 = count == count_max ? 10'h0 : _GEN_127; // @[PEArray.scala 202:32 PEArray.scala 203:15]
  wire [2:0] _GEN_331 = count == count_max ? 3'h0 : state; // @[PEArray.scala 202:32 PEArray.scala 204:15 PEArray.scala 100:22]
  wire [9:0] _GEN_865 = {{4'd0}, GRU_out_width}; // @[PEArray.scala 220:19]
  wire [9:0] _GEN_0 = count % _GEN_865; // @[PEArray.scala 220:19]
  wire [5:0] _T_36 = _GEN_0[5:0]; // @[PEArray.scala 220:19]
  wire [5:0] _T_38 = GRU_out_width - 6'h1; // @[PEArray.scala 220:55]
  wire [5:0] _GEN_334 = _T_36 == _T_38 ? _L0Index_T_2 : L0index_begin; // @[PEArray.scala 220:62 PEArray.scala 221:17 PEArray.scala 214:15]
  wire [5:0] _GEN_346 = _T_41 ? _GEN_334 : L0Index; // @[Conditional.scala 39:67 PEArray.scala 39:24]
  wire [9:0] _GEN_347 = _T_41 ? _GEN_330 : count; // @[Conditional.scala 39:67 PEArray.scala 101:22]
  wire [2:0] _GEN_348 = _T_41 ? _GEN_331 : state; // @[Conditional.scala 39:67 PEArray.scala 100:22]
  wire [5:0] _GEN_353 = _T_31 ? _GEN_334 : _GEN_346; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_354 = _T_31 ? _GEN_330 : _GEN_347; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_355 = _T_31 ? _GEN_331 : _GEN_348; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_356 = _T_22 ? _GEN_330 : _GEN_354; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_357 = _T_22 ? _GEN_329 : _GEN_353; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_458 = _T_22 ? _GEN_331 : _GEN_355; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_690 = _T_3 ? _GEN_118 : {{2'd0}, GRU_out_width}; // @[Conditional.scala 40:58 PEArray.scala 104:26]
  FP16MulAdder FP16MAC ( // @[PEArray.scala 72:23]
    .io_a(FP16MAC_io_a),
    .io_b(FP16MAC_io_b),
    .io_c(FP16MAC_io_c),
    .io_out(FP16MAC_io_out)
  );
  assign io_ToRightPE = mux3out_reg; // @[PEArray.scala 95:16]
  assign io_ToBelowPE = mux2out_reg; // @[PEArray.scala 94:16]
  assign FP16MAC_io_a = sel1 ? io_FromL1 : io_FromLeftPE; // @[PEArray.scala 50:14 PEArray.scala 50:23 PEArray.scala 51:24]
  assign FP16MAC_io_b = sel5 ? mux4out : _GEN_105; // @[PEArray.scala 77:13 PEArray.scala 78:18 PEArray.scala 81:18]
  assign FP16MAC_io_c = sel5 ? _GEN_105 : mux4out; // @[PEArray.scala 77:13 PEArray.scala 79:18 PEArray.scala 82:18]
  always @(posedge clock) begin
    if (reset) begin // @[PEArray.scala 39:24]
      L0Index <= 6'h0; // @[PEArray.scala 39:24]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h2; // @[PEArray.scala 159:15]
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h9; // @[PEArray.scala 181:15]
      end else begin
        L0Index <= _GEN_357;
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_0 <= _GEN_229;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_1 <= _GEN_230;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_2 <= _GEN_231;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_3 <= _GEN_232;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_4 <= _GEN_233;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_5 <= _GEN_234;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_6 <= _GEN_235;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_7 <= _GEN_236;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_8 <= _GEN_237;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_9 <= _GEN_238;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_10 <= _GEN_239;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_11 <= _GEN_240;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_12 <= _GEN_241;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_13 <= _GEN_242;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_14 <= _GEN_243;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_15 <= _GEN_244;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_16 <= _GEN_245;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_17 <= _GEN_246;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_18 <= _GEN_247;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_19 <= _GEN_248;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_20 <= _GEN_249;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_21 <= _GEN_250;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_22 <= _GEN_251;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_23 <= _GEN_252;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_24 <= _GEN_253;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_25 <= _GEN_254;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_26 <= _GEN_255;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_27 <= _GEN_256;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_28 <= _GEN_257;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_29 <= _GEN_258;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_30 <= _GEN_259;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_31 <= _GEN_260;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_32 <= _GEN_261;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_33 <= _GEN_262;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_34 <= _GEN_263;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_35 <= _GEN_264;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_36 <= _GEN_265;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_37 <= _GEN_266;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_38 <= _GEN_267;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_39 <= _GEN_268;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_40 <= _GEN_269;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_41 <= _GEN_270;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_42 <= _GEN_271;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_43 <= _GEN_272;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_44 <= _GEN_273;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_45 <= _GEN_274;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_46 <= _GEN_275;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_47 <= _GEN_276;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_48 <= _GEN_277;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_49 <= _GEN_278;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_50 <= _GEN_279;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_51 <= _GEN_280;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_52 <= _GEN_281;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_53 <= _GEN_282;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_54 <= _GEN_283;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_55 <= _GEN_284;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_56 <= _GEN_285;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_57 <= _GEN_286;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_58 <= _GEN_287;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_59 <= _GEN_288;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_60 <= _GEN_289;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_61 <= _GEN_290;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_62 <= _GEN_291;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_63 <= _GEN_292;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_64 <= _GEN_293;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_65 <= _GEN_294;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_66 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_67 <= _GEN_296;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_68 <= _GEN_297;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_69 <= _GEN_298;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_70 <= _GEN_299;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_71 <= _GEN_300;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_72 <= _GEN_301;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_73 <= _GEN_302;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_74 <= _GEN_303;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_75 <= _GEN_304;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_76 <= _GEN_305;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_77 <= _GEN_306;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_78 <= _GEN_307;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_79 <= _GEN_308;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_80 <= _GEN_309;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_81 <= _GEN_310;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_82 <= _GEN_311;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_83 <= _GEN_312;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_84 <= _GEN_313;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_85 <= _GEN_314;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_86 <= _GEN_315;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_87 <= _GEN_316;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_88 <= _GEN_317;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_89 <= _GEN_318;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_90 <= _GEN_319;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_91 <= _GEN_320;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_92 <= _GEN_321;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_93 <= _GEN_322;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_94 <= _GEN_323;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_95 <= _GEN_324;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_96 <= _GEN_325;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_97 <= _GEN_326;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_98 <= _GEN_327;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_99 <= _GEN_328;
          end
        end
      end
    end
    if (reset) begin // @[PEArray.scala 100:22]
      state <= 3'h0; // @[PEArray.scala 100:22]
    end else if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[5]) begin // @[PEArray.scala 116:57]
        if (_T_6) begin // @[Conditional.scala 40:58]
          state <= 3'h0; // @[PEArray.scala 120:19]
        end else begin
          state <= _GEN_113;
        end
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      if (count == 10'h33) begin // @[PEArray.scala 164:27]
        state <= 3'h0; // @[PEArray.scala 166:15]
      end
    end else if (_T_16) begin // @[Conditional.scala 39:67]
      state <= _GEN_126;
    end else begin
      state <= _GEN_458;
    end
    if (reset) begin // @[PEArray.scala 90:28]
      mux2out_reg <= 16'h0; // @[PEArray.scala 90:28]
    end else begin
      mux2out_reg <= MAC_out; // @[PEArray.scala 90:28]
    end
    if (reset) begin // @[PEArray.scala 91:28]
      mux3out_reg <= 16'h0; // @[PEArray.scala 91:28]
    end else if (sel3) begin // @[PEArray.scala 56:14]
      mux3out_reg <= MAC_out; // @[PEArray.scala 56:23]
    end else if (sel1) begin // @[PEArray.scala 50:14]
      mux3out_reg <= io_FromL1; // @[PEArray.scala 50:23]
    end else begin
      mux3out_reg <= io_FromLeftPE; // @[PEArray.scala 51:24]
    end
    if (reset) begin // @[PEArray.scala 101:22]
      count <= 10'h0; // @[PEArray.scala 101:22]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        if (count == 10'h33) begin // @[PEArray.scala 164:27]
          count <= 10'h0; // @[PEArray.scala 165:15]
        end else begin
          count <= _GEN_120;
        end
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        count <= _GEN_125;
      end else begin
        count <= _GEN_356;
      end
    end
    if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[5]) begin // @[PEArray.scala 116:57]
        count_max <= io_control_signal_count; // @[PEArray.scala 143:19]
      end
    end
    if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[5]) begin // @[PEArray.scala 116:57]
        L0index_begin <= io_control_signal_L0index; // @[PEArray.scala 144:23]
      end
    end
    GRU_out_width <= _GEN_690[5:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  L0Index = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  L0Memory_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  L0Memory_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  L0Memory_2 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  L0Memory_3 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  L0Memory_4 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  L0Memory_5 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  L0Memory_6 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  L0Memory_7 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  L0Memory_8 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  L0Memory_9 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  L0Memory_10 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  L0Memory_11 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  L0Memory_12 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  L0Memory_13 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  L0Memory_14 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  L0Memory_15 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  L0Memory_16 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  L0Memory_17 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  L0Memory_18 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  L0Memory_19 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  L0Memory_20 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  L0Memory_21 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  L0Memory_22 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  L0Memory_23 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  L0Memory_24 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  L0Memory_25 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  L0Memory_26 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  L0Memory_27 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  L0Memory_28 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  L0Memory_29 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  L0Memory_30 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  L0Memory_31 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  L0Memory_32 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  L0Memory_33 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  L0Memory_34 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  L0Memory_35 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  L0Memory_36 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  L0Memory_37 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  L0Memory_38 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  L0Memory_39 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  L0Memory_40 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  L0Memory_41 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  L0Memory_42 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  L0Memory_43 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  L0Memory_44 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  L0Memory_45 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  L0Memory_46 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  L0Memory_47 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  L0Memory_48 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  L0Memory_49 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  L0Memory_50 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  L0Memory_51 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  L0Memory_52 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  L0Memory_53 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  L0Memory_54 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  L0Memory_55 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  L0Memory_56 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  L0Memory_57 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  L0Memory_58 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  L0Memory_59 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  L0Memory_60 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  L0Memory_61 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  L0Memory_62 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  L0Memory_63 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  L0Memory_64 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  L0Memory_65 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  L0Memory_66 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  L0Memory_67 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  L0Memory_68 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  L0Memory_69 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  L0Memory_70 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  L0Memory_71 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  L0Memory_72 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  L0Memory_73 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  L0Memory_74 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  L0Memory_75 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  L0Memory_76 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  L0Memory_77 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  L0Memory_78 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  L0Memory_79 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  L0Memory_80 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  L0Memory_81 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  L0Memory_82 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  L0Memory_83 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  L0Memory_84 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  L0Memory_85 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  L0Memory_86 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  L0Memory_87 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  L0Memory_88 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  L0Memory_89 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  L0Memory_90 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  L0Memory_91 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  L0Memory_92 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  L0Memory_93 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  L0Memory_94 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  L0Memory_95 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  L0Memory_96 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  L0Memory_97 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  L0Memory_98 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  L0Memory_99 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  state = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  mux2out_reg = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  mux3out_reg = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  count = _RAND_104[9:0];
  _RAND_105 = {1{`RANDOM}};
  count_max = _RAND_105[9:0];
  _RAND_106 = {1{`RANDOM}};
  L0index_begin = _RAND_106[5:0];
  _RAND_107 = {1{`RANDOM}};
  GRU_out_width = _RAND_107[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PE_21(
  input         clock,
  input         reset,
  input  [15:0] io_FromAbovePE,
  input  [15:0] io_FromLeftPE,
  input  [15:0] io_FromL1,
  input  [11:0] io_control_signal_mask,
  output [15:0] io_ToRightPE,
  output [15:0] io_ToBelowPE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] FP16MAC_io_a; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_b; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_c; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_out; // @[PEArray.scala 72:23]
  reg [5:0] L0Index; // @[PEArray.scala 39:24]
  reg [15:0] L0Memory_0; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_1; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_2; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_3; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_4; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_5; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_6; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_7; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_8; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_9; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_10; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_11; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_12; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_13; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_14; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_15; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_16; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_17; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_18; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_19; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_20; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_21; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_22; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_23; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_24; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_25; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_26; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_27; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_28; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_29; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_30; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_31; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_32; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_33; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_34; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_35; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_36; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_37; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_38; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_39; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_40; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_41; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_42; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_43; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_44; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_45; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_46; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_47; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_48; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_49; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_50; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_51; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_52; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_53; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_54; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_55; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_56; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_57; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_58; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_59; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_60; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_61; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_62; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_63; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_64; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_65; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_66; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_67; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_68; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_69; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_70; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_71; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_72; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_73; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_74; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_75; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_76; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_77; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_78; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_79; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_80; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_81; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_82; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_83; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_84; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_85; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_86; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_87; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_88; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_89; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_90; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_91; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_92; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_93; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_94; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_95; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_96; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_97; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_98; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_99; // @[PEArray.scala 40:21]
  reg [2:0] state; // @[PEArray.scala 100:22]
  wire  _T_3 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_12 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_16 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_22 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_31 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_41 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_342 = _T_41 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 231:12 PEArray.scala 32:8]
  wire  _GEN_349 = _T_31 ? 1'h0 : _GEN_342; // @[Conditional.scala 39:67 PEArray.scala 208:12]
  wire  _GEN_459 = _T_22 | _GEN_349; // @[Conditional.scala 39:67 PEArray.scala 32:8]
  wire  _GEN_463 = _T_16 ? 1'h0 : _GEN_459; // @[Conditional.scala 39:67]
  wire  _GEN_572 = _T_12 | _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 149:12]
  wire  sel1 = _T_3 | _GEN_572; // @[Conditional.scala 40:58 PEArray.scala 108:12]
  wire [15:0] MAC_out = FP16MAC_io_out; // @[PEArray.scala 47:21 PEArray.scala 85:11]
  wire  _GEN_465 = _T_16 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 177:12]
  wire  _GEN_580 = _T_12 | _GEN_465; // @[Conditional.scala 39:67 PEArray.scala 34:8]
  wire  sel3 = _T_3 | _GEN_580; // @[Conditional.scala 40:58 PEArray.scala 110:12]
  wire [1:0] _GEN_344 = _T_41 ? 2'h2 : 2'h0; // @[Conditional.scala 39:67 PEArray.scala 233:12 PEArray.scala 35:8]
  wire [1:0] _GEN_351 = _T_31 ? 2'h2 : _GEN_344; // @[Conditional.scala 39:67 PEArray.scala 210:12]
  wire [1:0] _GEN_461 = _T_22 ? 2'h0 : _GEN_351; // @[Conditional.scala 39:67 PEArray.scala 35:8]
  wire [1:0] _GEN_466 = _T_16 ? 2'h0 : _GEN_461; // @[Conditional.scala 39:67 PEArray.scala 178:12]
  wire [1:0] _GEN_574 = _T_12 ? 2'h0 : _GEN_466; // @[Conditional.scala 39:67]
  wire [1:0] sel4 = _T_3 ? 2'h0 : _GEN_574; // @[Conditional.scala 40:58 PEArray.scala 111:12]
  wire [15:0] _GEN_3 = sel4 == 2'h2 ? io_FromL1 : 16'h0; // @[PEArray.scala 65:28 PEArray.scala 66:15 PEArray.scala 69:15]
  wire [15:0] _GEN_4 = sel4 == 2'h1 ? io_FromAbovePE : _GEN_3; // @[PEArray.scala 62:28 PEArray.scala 63:15]
  wire [15:0] mux4out = sel4 == 2'h0 ? 16'h0 : _GEN_4; // @[PEArray.scala 59:22 PEArray.scala 60:13]
  wire [15:0] _GEN_7 = 6'h1 == L0Index ? L0Memory_1 : L0Memory_0; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_8 = 6'h2 == L0Index ? L0Memory_2 : _GEN_7; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_9 = 6'h3 == L0Index ? L0Memory_3 : _GEN_8; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_10 = 6'h4 == L0Index ? L0Memory_4 : _GEN_9; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_11 = 6'h5 == L0Index ? L0Memory_5 : _GEN_10; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_12 = 6'h6 == L0Index ? L0Memory_6 : _GEN_11; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_13 = 6'h7 == L0Index ? L0Memory_7 : _GEN_12; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_14 = 6'h8 == L0Index ? L0Memory_8 : _GEN_13; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_15 = 6'h9 == L0Index ? L0Memory_9 : _GEN_14; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_16 = 6'ha == L0Index ? L0Memory_10 : _GEN_15; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_17 = 6'hb == L0Index ? L0Memory_11 : _GEN_16; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_18 = 6'hc == L0Index ? L0Memory_12 : _GEN_17; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_19 = 6'hd == L0Index ? L0Memory_13 : _GEN_18; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_20 = 6'he == L0Index ? L0Memory_14 : _GEN_19; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_21 = 6'hf == L0Index ? L0Memory_15 : _GEN_20; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_22 = 6'h10 == L0Index ? L0Memory_16 : _GEN_21; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_23 = 6'h11 == L0Index ? L0Memory_17 : _GEN_22; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_24 = 6'h12 == L0Index ? L0Memory_18 : _GEN_23; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_25 = 6'h13 == L0Index ? L0Memory_19 : _GEN_24; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_26 = 6'h14 == L0Index ? L0Memory_20 : _GEN_25; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_27 = 6'h15 == L0Index ? L0Memory_21 : _GEN_26; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_28 = 6'h16 == L0Index ? L0Memory_22 : _GEN_27; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_29 = 6'h17 == L0Index ? L0Memory_23 : _GEN_28; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_30 = 6'h18 == L0Index ? L0Memory_24 : _GEN_29; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_31 = 6'h19 == L0Index ? L0Memory_25 : _GEN_30; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_32 = 6'h1a == L0Index ? L0Memory_26 : _GEN_31; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_33 = 6'h1b == L0Index ? L0Memory_27 : _GEN_32; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_34 = 6'h1c == L0Index ? L0Memory_28 : _GEN_33; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_35 = 6'h1d == L0Index ? L0Memory_29 : _GEN_34; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_36 = 6'h1e == L0Index ? L0Memory_30 : _GEN_35; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_37 = 6'h1f == L0Index ? L0Memory_31 : _GEN_36; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_38 = 6'h20 == L0Index ? L0Memory_32 : _GEN_37; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_39 = 6'h21 == L0Index ? L0Memory_33 : _GEN_38; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_40 = 6'h22 == L0Index ? L0Memory_34 : _GEN_39; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_41 = 6'h23 == L0Index ? L0Memory_35 : _GEN_40; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_42 = 6'h24 == L0Index ? L0Memory_36 : _GEN_41; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_43 = 6'h25 == L0Index ? L0Memory_37 : _GEN_42; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_44 = 6'h26 == L0Index ? L0Memory_38 : _GEN_43; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_45 = 6'h27 == L0Index ? L0Memory_39 : _GEN_44; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_46 = 6'h28 == L0Index ? L0Memory_40 : _GEN_45; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_47 = 6'h29 == L0Index ? L0Memory_41 : _GEN_46; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_48 = 6'h2a == L0Index ? L0Memory_42 : _GEN_47; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_49 = 6'h2b == L0Index ? L0Memory_43 : _GEN_48; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_50 = 6'h2c == L0Index ? L0Memory_44 : _GEN_49; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_51 = 6'h2d == L0Index ? L0Memory_45 : _GEN_50; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_52 = 6'h2e == L0Index ? L0Memory_46 : _GEN_51; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_53 = 6'h2f == L0Index ? L0Memory_47 : _GEN_52; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_54 = 6'h30 == L0Index ? L0Memory_48 : _GEN_53; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_55 = 6'h31 == L0Index ? L0Memory_49 : _GEN_54; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_56 = 6'h32 == L0Index ? L0Memory_50 : _GEN_55; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_57 = 6'h33 == L0Index ? L0Memory_51 : _GEN_56; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_58 = 6'h34 == L0Index ? L0Memory_52 : _GEN_57; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_59 = 6'h35 == L0Index ? L0Memory_53 : _GEN_58; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_60 = 6'h36 == L0Index ? L0Memory_54 : _GEN_59; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_61 = 6'h37 == L0Index ? L0Memory_55 : _GEN_60; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_62 = 6'h38 == L0Index ? L0Memory_56 : _GEN_61; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_63 = 6'h39 == L0Index ? L0Memory_57 : _GEN_62; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_64 = 6'h3a == L0Index ? L0Memory_58 : _GEN_63; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_65 = 6'h3b == L0Index ? L0Memory_59 : _GEN_64; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_66 = 6'h3c == L0Index ? L0Memory_60 : _GEN_65; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_67 = 6'h3d == L0Index ? L0Memory_61 : _GEN_66; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_68 = 6'h3e == L0Index ? L0Memory_62 : _GEN_67; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_69 = 6'h3f == L0Index ? L0Memory_63 : _GEN_68; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [6:0] _GEN_793 = {{1'd0}, L0Index}; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_70 = 7'h40 == _GEN_793 ? L0Memory_64 : _GEN_69; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_71 = 7'h41 == _GEN_793 ? L0Memory_65 : _GEN_70; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_72 = 7'h42 == _GEN_793 ? L0Memory_66 : _GEN_71; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_73 = 7'h43 == _GEN_793 ? L0Memory_67 : _GEN_72; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_74 = 7'h44 == _GEN_793 ? L0Memory_68 : _GEN_73; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_75 = 7'h45 == _GEN_793 ? L0Memory_69 : _GEN_74; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_76 = 7'h46 == _GEN_793 ? L0Memory_70 : _GEN_75; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_77 = 7'h47 == _GEN_793 ? L0Memory_71 : _GEN_76; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_78 = 7'h48 == _GEN_793 ? L0Memory_72 : _GEN_77; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_79 = 7'h49 == _GEN_793 ? L0Memory_73 : _GEN_78; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_80 = 7'h4a == _GEN_793 ? L0Memory_74 : _GEN_79; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_81 = 7'h4b == _GEN_793 ? L0Memory_75 : _GEN_80; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_82 = 7'h4c == _GEN_793 ? L0Memory_76 : _GEN_81; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_83 = 7'h4d == _GEN_793 ? L0Memory_77 : _GEN_82; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_84 = 7'h4e == _GEN_793 ? L0Memory_78 : _GEN_83; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_85 = 7'h4f == _GEN_793 ? L0Memory_79 : _GEN_84; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_86 = 7'h50 == _GEN_793 ? L0Memory_80 : _GEN_85; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_87 = 7'h51 == _GEN_793 ? L0Memory_81 : _GEN_86; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_88 = 7'h52 == _GEN_793 ? L0Memory_82 : _GEN_87; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_89 = 7'h53 == _GEN_793 ? L0Memory_83 : _GEN_88; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_90 = 7'h54 == _GEN_793 ? L0Memory_84 : _GEN_89; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_91 = 7'h55 == _GEN_793 ? L0Memory_85 : _GEN_90; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_92 = 7'h56 == _GEN_793 ? L0Memory_86 : _GEN_91; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_93 = 7'h57 == _GEN_793 ? L0Memory_87 : _GEN_92; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_94 = 7'h58 == _GEN_793 ? L0Memory_88 : _GEN_93; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_95 = 7'h59 == _GEN_793 ? L0Memory_89 : _GEN_94; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_96 = 7'h5a == _GEN_793 ? L0Memory_90 : _GEN_95; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_97 = 7'h5b == _GEN_793 ? L0Memory_91 : _GEN_96; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_98 = 7'h5c == _GEN_793 ? L0Memory_92 : _GEN_97; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_99 = 7'h5d == _GEN_793 ? L0Memory_93 : _GEN_98; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_100 = 7'h5e == _GEN_793 ? L0Memory_94 : _GEN_99; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_101 = 7'h5f == _GEN_793 ? L0Memory_95 : _GEN_100; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_102 = 7'h60 == _GEN_793 ? L0Memory_96 : _GEN_101; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_103 = 7'h61 == _GEN_793 ? L0Memory_97 : _GEN_102; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_104 = 7'h62 == _GEN_793 ? L0Memory_98 : _GEN_103; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_105 = 7'h63 == _GEN_793 ? L0Memory_99 : _GEN_104; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire  _GEN_575 = _T_12 ? 1'h0 : _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 157:12]
  wire  sel5 = _T_3 ? 1'h0 : _GEN_575; // @[Conditional.scala 40:58 PEArray.scala 112:12]
  reg [15:0] mux2out_reg; // @[PEArray.scala 90:28]
  reg [15:0] mux3out_reg; // @[PEArray.scala 91:28]
  reg [9:0] count; // @[PEArray.scala 101:22]
  reg [5:0] GRU_out_width; // @[PEArray.scala 104:26]
  wire [7:0] _GEN_118 = io_control_signal_mask[4] ? 8'h0 : {{2'd0}, GRU_out_width}; // @[PEArray.scala 116:57 PEArray.scala 145:23 PEArray.scala 104:26]
  wire [9:0] _count_T_1 = count + 10'h1; // @[PEArray.scala 162:24]
  wire [9:0] _GEN_120 = count != 10'h33 ? _count_T_1 : count; // @[PEArray.scala 161:27 PEArray.scala 162:15 PEArray.scala 101:22]
  wire [9:0] _GEN_124 = count != 10'h188 ? _count_T_1 : count; // @[PEArray.scala 183:28 PEArray.scala 184:15 PEArray.scala 101:22]
  wire [9:0] _GEN_125 = count == 10'h188 ? 10'h0 : _GEN_124; // @[PEArray.scala 186:28 PEArray.scala 187:15]
  wire [2:0] _GEN_126 = count == 10'h188 ? 3'h0 : state; // @[PEArray.scala 186:28 PEArray.scala 188:15 PEArray.scala 100:22]
  wire [9:0] _GEN_127 = count != 10'h0 ? _count_T_1 : count; // @[PEArray.scala 192:32 PEArray.scala 193:15 PEArray.scala 101:22]
  wire  _T_24 = count == 10'h0; // @[PEArray.scala 195:18]
  wire [5:0] _GEN_128 = count == 10'h0 ? 6'h0 : L0Index; // @[PEArray.scala 195:26 PEArray.scala 196:17 PEArray.scala 39:24]
  wire [9:0] _T_27 = 10'h0 - 10'h1; // @[PEArray.scala 198:51]
  wire [15:0] _GEN_129 = 6'h0 == L0Index ? io_FromL1 : L0Memory_0; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_130 = 6'h1 == L0Index ? io_FromL1 : L0Memory_1; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_131 = 6'h2 == L0Index ? io_FromL1 : L0Memory_2; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_132 = 6'h3 == L0Index ? io_FromL1 : L0Memory_3; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_133 = 6'h4 == L0Index ? io_FromL1 : L0Memory_4; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_134 = 6'h5 == L0Index ? io_FromL1 : L0Memory_5; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_135 = 6'h6 == L0Index ? io_FromL1 : L0Memory_6; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_136 = 6'h7 == L0Index ? io_FromL1 : L0Memory_7; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_137 = 6'h8 == L0Index ? io_FromL1 : L0Memory_8; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_138 = 6'h9 == L0Index ? io_FromL1 : L0Memory_9; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_139 = 6'ha == L0Index ? io_FromL1 : L0Memory_10; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_140 = 6'hb == L0Index ? io_FromL1 : L0Memory_11; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_141 = 6'hc == L0Index ? io_FromL1 : L0Memory_12; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_142 = 6'hd == L0Index ? io_FromL1 : L0Memory_13; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_143 = 6'he == L0Index ? io_FromL1 : L0Memory_14; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_144 = 6'hf == L0Index ? io_FromL1 : L0Memory_15; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_145 = 6'h10 == L0Index ? io_FromL1 : L0Memory_16; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_146 = 6'h11 == L0Index ? io_FromL1 : L0Memory_17; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_147 = 6'h12 == L0Index ? io_FromL1 : L0Memory_18; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_148 = 6'h13 == L0Index ? io_FromL1 : L0Memory_19; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_149 = 6'h14 == L0Index ? io_FromL1 : L0Memory_20; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_150 = 6'h15 == L0Index ? io_FromL1 : L0Memory_21; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_151 = 6'h16 == L0Index ? io_FromL1 : L0Memory_22; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_152 = 6'h17 == L0Index ? io_FromL1 : L0Memory_23; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_153 = 6'h18 == L0Index ? io_FromL1 : L0Memory_24; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_154 = 6'h19 == L0Index ? io_FromL1 : L0Memory_25; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_155 = 6'h1a == L0Index ? io_FromL1 : L0Memory_26; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_156 = 6'h1b == L0Index ? io_FromL1 : L0Memory_27; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_157 = 6'h1c == L0Index ? io_FromL1 : L0Memory_28; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_158 = 6'h1d == L0Index ? io_FromL1 : L0Memory_29; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_159 = 6'h1e == L0Index ? io_FromL1 : L0Memory_30; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_160 = 6'h1f == L0Index ? io_FromL1 : L0Memory_31; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_161 = 6'h20 == L0Index ? io_FromL1 : L0Memory_32; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_162 = 6'h21 == L0Index ? io_FromL1 : L0Memory_33; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_163 = 6'h22 == L0Index ? io_FromL1 : L0Memory_34; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_164 = 6'h23 == L0Index ? io_FromL1 : L0Memory_35; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_165 = 6'h24 == L0Index ? io_FromL1 : L0Memory_36; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_166 = 6'h25 == L0Index ? io_FromL1 : L0Memory_37; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_167 = 6'h26 == L0Index ? io_FromL1 : L0Memory_38; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_168 = 6'h27 == L0Index ? io_FromL1 : L0Memory_39; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_169 = 6'h28 == L0Index ? io_FromL1 : L0Memory_40; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_170 = 6'h29 == L0Index ? io_FromL1 : L0Memory_41; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_171 = 6'h2a == L0Index ? io_FromL1 : L0Memory_42; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_172 = 6'h2b == L0Index ? io_FromL1 : L0Memory_43; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_173 = 6'h2c == L0Index ? io_FromL1 : L0Memory_44; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_174 = 6'h2d == L0Index ? io_FromL1 : L0Memory_45; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_175 = 6'h2e == L0Index ? io_FromL1 : L0Memory_46; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_176 = 6'h2f == L0Index ? io_FromL1 : L0Memory_47; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_177 = 6'h30 == L0Index ? io_FromL1 : L0Memory_48; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_178 = 6'h31 == L0Index ? io_FromL1 : L0Memory_49; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_179 = 6'h32 == L0Index ? io_FromL1 : L0Memory_50; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_180 = 6'h33 == L0Index ? io_FromL1 : L0Memory_51; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_181 = 6'h34 == L0Index ? io_FromL1 : L0Memory_52; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_182 = 6'h35 == L0Index ? io_FromL1 : L0Memory_53; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_183 = 6'h36 == L0Index ? io_FromL1 : L0Memory_54; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_184 = 6'h37 == L0Index ? io_FromL1 : L0Memory_55; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_185 = 6'h38 == L0Index ? io_FromL1 : L0Memory_56; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_186 = 6'h39 == L0Index ? io_FromL1 : L0Memory_57; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_187 = 6'h3a == L0Index ? io_FromL1 : L0Memory_58; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_188 = 6'h3b == L0Index ? io_FromL1 : L0Memory_59; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_189 = 6'h3c == L0Index ? io_FromL1 : L0Memory_60; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_190 = 6'h3d == L0Index ? io_FromL1 : L0Memory_61; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_191 = 6'h3e == L0Index ? io_FromL1 : L0Memory_62; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_192 = 6'h3f == L0Index ? io_FromL1 : L0Memory_63; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_193 = 7'h40 == _GEN_793 ? io_FromL1 : L0Memory_64; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_194 = 7'h41 == _GEN_793 ? io_FromL1 : L0Memory_65; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_195 = 7'h42 == _GEN_793 ? io_FromL1 : L0Memory_66; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_196 = 7'h43 == _GEN_793 ? io_FromL1 : L0Memory_67; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_197 = 7'h44 == _GEN_793 ? io_FromL1 : L0Memory_68; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_198 = 7'h45 == _GEN_793 ? io_FromL1 : L0Memory_69; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_199 = 7'h46 == _GEN_793 ? io_FromL1 : L0Memory_70; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_200 = 7'h47 == _GEN_793 ? io_FromL1 : L0Memory_71; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_201 = 7'h48 == _GEN_793 ? io_FromL1 : L0Memory_72; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_202 = 7'h49 == _GEN_793 ? io_FromL1 : L0Memory_73; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_203 = 7'h4a == _GEN_793 ? io_FromL1 : L0Memory_74; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_204 = 7'h4b == _GEN_793 ? io_FromL1 : L0Memory_75; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_205 = 7'h4c == _GEN_793 ? io_FromL1 : L0Memory_76; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_206 = 7'h4d == _GEN_793 ? io_FromL1 : L0Memory_77; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_207 = 7'h4e == _GEN_793 ? io_FromL1 : L0Memory_78; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_208 = 7'h4f == _GEN_793 ? io_FromL1 : L0Memory_79; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_209 = 7'h50 == _GEN_793 ? io_FromL1 : L0Memory_80; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_210 = 7'h51 == _GEN_793 ? io_FromL1 : L0Memory_81; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_211 = 7'h52 == _GEN_793 ? io_FromL1 : L0Memory_82; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_212 = 7'h53 == _GEN_793 ? io_FromL1 : L0Memory_83; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_213 = 7'h54 == _GEN_793 ? io_FromL1 : L0Memory_84; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_214 = 7'h55 == _GEN_793 ? io_FromL1 : L0Memory_85; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_215 = 7'h56 == _GEN_793 ? io_FromL1 : L0Memory_86; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_216 = 7'h57 == _GEN_793 ? io_FromL1 : L0Memory_87; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_217 = 7'h58 == _GEN_793 ? io_FromL1 : L0Memory_88; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_218 = 7'h59 == _GEN_793 ? io_FromL1 : L0Memory_89; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_219 = 7'h5a == _GEN_793 ? io_FromL1 : L0Memory_90; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_220 = 7'h5b == _GEN_793 ? io_FromL1 : L0Memory_91; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_221 = 7'h5c == _GEN_793 ? io_FromL1 : L0Memory_92; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_222 = 7'h5d == _GEN_793 ? io_FromL1 : L0Memory_93; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_223 = 7'h5e == _GEN_793 ? io_FromL1 : L0Memory_94; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_224 = 7'h5f == _GEN_793 ? io_FromL1 : L0Memory_95; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_225 = 7'h60 == _GEN_793 ? io_FromL1 : L0Memory_96; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_226 = 7'h61 == _GEN_793 ? io_FromL1 : L0Memory_97; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_227 = 7'h62 == _GEN_793 ? io_FromL1 : L0Memory_98; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_228 = 7'h63 == _GEN_793 ? io_FromL1 : L0Memory_99; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [5:0] _L0Index_T_2 = L0Index + 6'h1; // @[PEArray.scala 200:28]
  wire [15:0] _GEN_229 = count >= 10'h1 & count <= _T_27 ? _GEN_129 : L0Memory_0; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_230 = count >= 10'h1 & count <= _T_27 ? _GEN_130 : L0Memory_1; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_231 = count >= 10'h1 & count <= _T_27 ? _GEN_131 : L0Memory_2; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_232 = count >= 10'h1 & count <= _T_27 ? _GEN_132 : L0Memory_3; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_233 = count >= 10'h1 & count <= _T_27 ? _GEN_133 : L0Memory_4; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_234 = count >= 10'h1 & count <= _T_27 ? _GEN_134 : L0Memory_5; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_235 = count >= 10'h1 & count <= _T_27 ? _GEN_135 : L0Memory_6; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_236 = count >= 10'h1 & count <= _T_27 ? _GEN_136 : L0Memory_7; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_237 = count >= 10'h1 & count <= _T_27 ? _GEN_137 : L0Memory_8; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_238 = count >= 10'h1 & count <= _T_27 ? _GEN_138 : L0Memory_9; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_239 = count >= 10'h1 & count <= _T_27 ? _GEN_139 : L0Memory_10; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_240 = count >= 10'h1 & count <= _T_27 ? _GEN_140 : L0Memory_11; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_241 = count >= 10'h1 & count <= _T_27 ? _GEN_141 : L0Memory_12; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_242 = count >= 10'h1 & count <= _T_27 ? _GEN_142 : L0Memory_13; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_243 = count >= 10'h1 & count <= _T_27 ? _GEN_143 : L0Memory_14; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_244 = count >= 10'h1 & count <= _T_27 ? _GEN_144 : L0Memory_15; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_245 = count >= 10'h1 & count <= _T_27 ? _GEN_145 : L0Memory_16; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_246 = count >= 10'h1 & count <= _T_27 ? _GEN_146 : L0Memory_17; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_247 = count >= 10'h1 & count <= _T_27 ? _GEN_147 : L0Memory_18; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_248 = count >= 10'h1 & count <= _T_27 ? _GEN_148 : L0Memory_19; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_249 = count >= 10'h1 & count <= _T_27 ? _GEN_149 : L0Memory_20; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_250 = count >= 10'h1 & count <= _T_27 ? _GEN_150 : L0Memory_21; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_251 = count >= 10'h1 & count <= _T_27 ? _GEN_151 : L0Memory_22; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_252 = count >= 10'h1 & count <= _T_27 ? _GEN_152 : L0Memory_23; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_253 = count >= 10'h1 & count <= _T_27 ? _GEN_153 : L0Memory_24; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_254 = count >= 10'h1 & count <= _T_27 ? _GEN_154 : L0Memory_25; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_255 = count >= 10'h1 & count <= _T_27 ? _GEN_155 : L0Memory_26; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_256 = count >= 10'h1 & count <= _T_27 ? _GEN_156 : L0Memory_27; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_257 = count >= 10'h1 & count <= _T_27 ? _GEN_157 : L0Memory_28; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_258 = count >= 10'h1 & count <= _T_27 ? _GEN_158 : L0Memory_29; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_259 = count >= 10'h1 & count <= _T_27 ? _GEN_159 : L0Memory_30; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_260 = count >= 10'h1 & count <= _T_27 ? _GEN_160 : L0Memory_31; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_261 = count >= 10'h1 & count <= _T_27 ? _GEN_161 : L0Memory_32; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_262 = count >= 10'h1 & count <= _T_27 ? _GEN_162 : L0Memory_33; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_263 = count >= 10'h1 & count <= _T_27 ? _GEN_163 : L0Memory_34; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_264 = count >= 10'h1 & count <= _T_27 ? _GEN_164 : L0Memory_35; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_265 = count >= 10'h1 & count <= _T_27 ? _GEN_165 : L0Memory_36; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_266 = count >= 10'h1 & count <= _T_27 ? _GEN_166 : L0Memory_37; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_267 = count >= 10'h1 & count <= _T_27 ? _GEN_167 : L0Memory_38; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_268 = count >= 10'h1 & count <= _T_27 ? _GEN_168 : L0Memory_39; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_269 = count >= 10'h1 & count <= _T_27 ? _GEN_169 : L0Memory_40; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_270 = count >= 10'h1 & count <= _T_27 ? _GEN_170 : L0Memory_41; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_271 = count >= 10'h1 & count <= _T_27 ? _GEN_171 : L0Memory_42; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_272 = count >= 10'h1 & count <= _T_27 ? _GEN_172 : L0Memory_43; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_273 = count >= 10'h1 & count <= _T_27 ? _GEN_173 : L0Memory_44; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_274 = count >= 10'h1 & count <= _T_27 ? _GEN_174 : L0Memory_45; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_275 = count >= 10'h1 & count <= _T_27 ? _GEN_175 : L0Memory_46; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_276 = count >= 10'h1 & count <= _T_27 ? _GEN_176 : L0Memory_47; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_277 = count >= 10'h1 & count <= _T_27 ? _GEN_177 : L0Memory_48; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_278 = count >= 10'h1 & count <= _T_27 ? _GEN_178 : L0Memory_49; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_279 = count >= 10'h1 & count <= _T_27 ? _GEN_179 : L0Memory_50; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_280 = count >= 10'h1 & count <= _T_27 ? _GEN_180 : L0Memory_51; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_281 = count >= 10'h1 & count <= _T_27 ? _GEN_181 : L0Memory_52; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_282 = count >= 10'h1 & count <= _T_27 ? _GEN_182 : L0Memory_53; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_283 = count >= 10'h1 & count <= _T_27 ? _GEN_183 : L0Memory_54; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_284 = count >= 10'h1 & count <= _T_27 ? _GEN_184 : L0Memory_55; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_285 = count >= 10'h1 & count <= _T_27 ? _GEN_185 : L0Memory_56; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_286 = count >= 10'h1 & count <= _T_27 ? _GEN_186 : L0Memory_57; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_287 = count >= 10'h1 & count <= _T_27 ? _GEN_187 : L0Memory_58; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_288 = count >= 10'h1 & count <= _T_27 ? _GEN_188 : L0Memory_59; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_289 = count >= 10'h1 & count <= _T_27 ? _GEN_189 : L0Memory_60; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_290 = count >= 10'h1 & count <= _T_27 ? _GEN_190 : L0Memory_61; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_291 = count >= 10'h1 & count <= _T_27 ? _GEN_191 : L0Memory_62; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_292 = count >= 10'h1 & count <= _T_27 ? _GEN_192 : L0Memory_63; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_293 = count >= 10'h1 & count <= _T_27 ? _GEN_193 : L0Memory_64; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_294 = count >= 10'h1 & count <= _T_27 ? _GEN_194 : L0Memory_65; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_295 = count >= 10'h1 & count <= _T_27 ? _GEN_195 : L0Memory_66; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_296 = count >= 10'h1 & count <= _T_27 ? _GEN_196 : L0Memory_67; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_297 = count >= 10'h1 & count <= _T_27 ? _GEN_197 : L0Memory_68; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_298 = count >= 10'h1 & count <= _T_27 ? _GEN_198 : L0Memory_69; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_299 = count >= 10'h1 & count <= _T_27 ? _GEN_199 : L0Memory_70; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_300 = count >= 10'h1 & count <= _T_27 ? _GEN_200 : L0Memory_71; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_301 = count >= 10'h1 & count <= _T_27 ? _GEN_201 : L0Memory_72; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_302 = count >= 10'h1 & count <= _T_27 ? _GEN_202 : L0Memory_73; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_303 = count >= 10'h1 & count <= _T_27 ? _GEN_203 : L0Memory_74; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_304 = count >= 10'h1 & count <= _T_27 ? _GEN_204 : L0Memory_75; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_305 = count >= 10'h1 & count <= _T_27 ? _GEN_205 : L0Memory_76; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_306 = count >= 10'h1 & count <= _T_27 ? _GEN_206 : L0Memory_77; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_307 = count >= 10'h1 & count <= _T_27 ? _GEN_207 : L0Memory_78; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_308 = count >= 10'h1 & count <= _T_27 ? _GEN_208 : L0Memory_79; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_309 = count >= 10'h1 & count <= _T_27 ? _GEN_209 : L0Memory_80; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_310 = count >= 10'h1 & count <= _T_27 ? _GEN_210 : L0Memory_81; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_311 = count >= 10'h1 & count <= _T_27 ? _GEN_211 : L0Memory_82; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_312 = count >= 10'h1 & count <= _T_27 ? _GEN_212 : L0Memory_83; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_313 = count >= 10'h1 & count <= _T_27 ? _GEN_213 : L0Memory_84; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_314 = count >= 10'h1 & count <= _T_27 ? _GEN_214 : L0Memory_85; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_315 = count >= 10'h1 & count <= _T_27 ? _GEN_215 : L0Memory_86; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_316 = count >= 10'h1 & count <= _T_27 ? _GEN_216 : L0Memory_87; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_317 = count >= 10'h1 & count <= _T_27 ? _GEN_217 : L0Memory_88; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_318 = count >= 10'h1 & count <= _T_27 ? _GEN_218 : L0Memory_89; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_319 = count >= 10'h1 & count <= _T_27 ? _GEN_219 : L0Memory_90; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_320 = count >= 10'h1 & count <= _T_27 ? _GEN_220 : L0Memory_91; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_321 = count >= 10'h1 & count <= _T_27 ? _GEN_221 : L0Memory_92; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_322 = count >= 10'h1 & count <= _T_27 ? _GEN_222 : L0Memory_93; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_323 = count >= 10'h1 & count <= _T_27 ? _GEN_223 : L0Memory_94; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_324 = count >= 10'h1 & count <= _T_27 ? _GEN_224 : L0Memory_95; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_325 = count >= 10'h1 & count <= _T_27 ? _GEN_225 : L0Memory_96; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_326 = count >= 10'h1 & count <= _T_27 ? _GEN_226 : L0Memory_97; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_327 = count >= 10'h1 & count <= _T_27 ? _GEN_227 : L0Memory_98; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_328 = count >= 10'h1 & count <= _T_27 ? _GEN_228 : L0Memory_99; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [5:0] _GEN_329 = count >= 10'h1 & count <= _T_27 ? _L0Index_T_2 : _GEN_128; // @[PEArray.scala 198:59 PEArray.scala 200:17]
  wire [9:0] _GEN_330 = _T_24 ? 10'h0 : _GEN_127; // @[PEArray.scala 202:32 PEArray.scala 203:15]
  wire [2:0] _GEN_331 = _T_24 ? 3'h0 : state; // @[PEArray.scala 202:32 PEArray.scala 204:15 PEArray.scala 100:22]
  wire [9:0] _GEN_865 = {{4'd0}, GRU_out_width}; // @[PEArray.scala 220:19]
  wire [9:0] _GEN_0 = count % _GEN_865; // @[PEArray.scala 220:19]
  wire [5:0] _T_36 = _GEN_0[5:0]; // @[PEArray.scala 220:19]
  wire [5:0] _T_38 = GRU_out_width - 6'h1; // @[PEArray.scala 220:55]
  wire [5:0] _GEN_334 = _T_36 == _T_38 ? _L0Index_T_2 : 6'h0; // @[PEArray.scala 220:62 PEArray.scala 221:17 PEArray.scala 214:15]
  wire [5:0] _GEN_346 = _T_41 ? _GEN_334 : L0Index; // @[Conditional.scala 39:67 PEArray.scala 39:24]
  wire [9:0] _GEN_347 = _T_41 ? _GEN_330 : count; // @[Conditional.scala 39:67 PEArray.scala 101:22]
  wire [2:0] _GEN_348 = _T_41 ? _GEN_331 : state; // @[Conditional.scala 39:67 PEArray.scala 100:22]
  wire [5:0] _GEN_353 = _T_31 ? _GEN_334 : _GEN_346; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_354 = _T_31 ? _GEN_330 : _GEN_347; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_355 = _T_31 ? _GEN_331 : _GEN_348; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_356 = _T_22 ? _GEN_330 : _GEN_354; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_357 = _T_22 ? _GEN_329 : _GEN_353; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_458 = _T_22 ? _GEN_331 : _GEN_355; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_690 = _T_3 ? _GEN_118 : {{2'd0}, GRU_out_width}; // @[Conditional.scala 40:58 PEArray.scala 104:26]
  FP16MulAdder FP16MAC ( // @[PEArray.scala 72:23]
    .io_a(FP16MAC_io_a),
    .io_b(FP16MAC_io_b),
    .io_c(FP16MAC_io_c),
    .io_out(FP16MAC_io_out)
  );
  assign io_ToRightPE = mux3out_reg; // @[PEArray.scala 95:16]
  assign io_ToBelowPE = mux2out_reg; // @[PEArray.scala 94:16]
  assign FP16MAC_io_a = sel1 ? io_FromL1 : io_FromLeftPE; // @[PEArray.scala 50:14 PEArray.scala 50:23 PEArray.scala 51:24]
  assign FP16MAC_io_b = sel5 ? mux4out : _GEN_105; // @[PEArray.scala 77:13 PEArray.scala 78:18 PEArray.scala 81:18]
  assign FP16MAC_io_c = sel5 ? _GEN_105 : mux4out; // @[PEArray.scala 77:13 PEArray.scala 79:18 PEArray.scala 82:18]
  always @(posedge clock) begin
    if (reset) begin // @[PEArray.scala 39:24]
      L0Index <= 6'h0; // @[PEArray.scala 39:24]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h0; // @[PEArray.scala 159:15]
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        L0Index <= 6'ha; // @[PEArray.scala 181:15]
      end else begin
        L0Index <= _GEN_357;
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_0 <= _GEN_229;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_1 <= _GEN_230;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_2 <= _GEN_231;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_3 <= _GEN_232;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_4 <= _GEN_233;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_5 <= _GEN_234;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_6 <= _GEN_235;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_7 <= _GEN_236;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_8 <= _GEN_237;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_9 <= _GEN_238;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_10 <= _GEN_239;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_11 <= _GEN_240;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_12 <= _GEN_241;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_13 <= _GEN_242;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_14 <= _GEN_243;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_15 <= _GEN_244;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_16 <= _GEN_245;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_17 <= _GEN_246;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_18 <= _GEN_247;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_19 <= _GEN_248;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_20 <= _GEN_249;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_21 <= _GEN_250;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_22 <= _GEN_251;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_23 <= _GEN_252;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_24 <= _GEN_253;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_25 <= _GEN_254;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_26 <= _GEN_255;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_27 <= _GEN_256;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_28 <= _GEN_257;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_29 <= _GEN_258;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_30 <= _GEN_259;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_31 <= _GEN_260;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_32 <= _GEN_261;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_33 <= _GEN_262;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_34 <= _GEN_263;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_35 <= _GEN_264;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_36 <= _GEN_265;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_37 <= _GEN_266;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_38 <= _GEN_267;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_39 <= _GEN_268;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_40 <= _GEN_269;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_41 <= _GEN_270;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_42 <= _GEN_271;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_43 <= _GEN_272;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_44 <= _GEN_273;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_45 <= _GEN_274;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_46 <= _GEN_275;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_47 <= _GEN_276;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_48 <= _GEN_277;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_49 <= _GEN_278;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_50 <= _GEN_279;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_51 <= _GEN_280;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_52 <= _GEN_281;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_53 <= _GEN_282;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_54 <= _GEN_283;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_55 <= _GEN_284;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_56 <= _GEN_285;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_57 <= _GEN_286;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_58 <= _GEN_287;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_59 <= _GEN_288;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_60 <= _GEN_289;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_61 <= _GEN_290;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_62 <= _GEN_291;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_63 <= _GEN_292;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_64 <= _GEN_293;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_65 <= _GEN_294;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_66 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_67 <= _GEN_296;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_68 <= _GEN_297;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_69 <= _GEN_298;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_70 <= _GEN_299;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_71 <= _GEN_300;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_72 <= _GEN_301;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_73 <= _GEN_302;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_74 <= _GEN_303;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_75 <= _GEN_304;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_76 <= _GEN_305;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_77 <= _GEN_306;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_78 <= _GEN_307;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_79 <= _GEN_308;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_80 <= _GEN_309;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_81 <= _GEN_310;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_82 <= _GEN_311;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_83 <= _GEN_312;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_84 <= _GEN_313;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_85 <= _GEN_314;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_86 <= _GEN_315;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_87 <= _GEN_316;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_88 <= _GEN_317;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_89 <= _GEN_318;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_90 <= _GEN_319;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_91 <= _GEN_320;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_92 <= _GEN_321;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_93 <= _GEN_322;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_94 <= _GEN_323;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_95 <= _GEN_324;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_96 <= _GEN_325;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_97 <= _GEN_326;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_98 <= _GEN_327;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_99 <= _GEN_328;
          end
        end
      end
    end
    if (reset) begin // @[PEArray.scala 100:22]
      state <= 3'h0; // @[PEArray.scala 100:22]
    end else if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[4]) begin // @[PEArray.scala 116:57]
        state <= 3'h1;
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      if (count == 10'h33) begin // @[PEArray.scala 164:27]
        state <= 3'h0; // @[PEArray.scala 166:15]
      end
    end else if (_T_16) begin // @[Conditional.scala 39:67]
      state <= _GEN_126;
    end else begin
      state <= _GEN_458;
    end
    if (reset) begin // @[PEArray.scala 90:28]
      mux2out_reg <= 16'h0; // @[PEArray.scala 90:28]
    end else begin
      mux2out_reg <= MAC_out; // @[PEArray.scala 90:28]
    end
    if (reset) begin // @[PEArray.scala 91:28]
      mux3out_reg <= 16'h0; // @[PEArray.scala 91:28]
    end else if (sel3) begin // @[PEArray.scala 56:14]
      mux3out_reg <= MAC_out; // @[PEArray.scala 56:23]
    end else if (sel1) begin // @[PEArray.scala 50:14]
      mux3out_reg <= io_FromL1; // @[PEArray.scala 50:23]
    end else begin
      mux3out_reg <= io_FromLeftPE; // @[PEArray.scala 51:24]
    end
    if (reset) begin // @[PEArray.scala 101:22]
      count <= 10'h0; // @[PEArray.scala 101:22]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        if (count == 10'h33) begin // @[PEArray.scala 164:27]
          count <= 10'h0; // @[PEArray.scala 165:15]
        end else begin
          count <= _GEN_120;
        end
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        count <= _GEN_125;
      end else begin
        count <= _GEN_356;
      end
    end
    GRU_out_width <= _GEN_690[5:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  L0Index = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  L0Memory_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  L0Memory_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  L0Memory_2 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  L0Memory_3 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  L0Memory_4 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  L0Memory_5 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  L0Memory_6 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  L0Memory_7 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  L0Memory_8 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  L0Memory_9 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  L0Memory_10 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  L0Memory_11 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  L0Memory_12 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  L0Memory_13 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  L0Memory_14 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  L0Memory_15 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  L0Memory_16 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  L0Memory_17 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  L0Memory_18 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  L0Memory_19 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  L0Memory_20 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  L0Memory_21 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  L0Memory_22 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  L0Memory_23 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  L0Memory_24 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  L0Memory_25 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  L0Memory_26 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  L0Memory_27 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  L0Memory_28 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  L0Memory_29 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  L0Memory_30 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  L0Memory_31 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  L0Memory_32 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  L0Memory_33 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  L0Memory_34 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  L0Memory_35 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  L0Memory_36 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  L0Memory_37 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  L0Memory_38 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  L0Memory_39 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  L0Memory_40 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  L0Memory_41 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  L0Memory_42 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  L0Memory_43 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  L0Memory_44 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  L0Memory_45 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  L0Memory_46 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  L0Memory_47 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  L0Memory_48 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  L0Memory_49 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  L0Memory_50 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  L0Memory_51 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  L0Memory_52 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  L0Memory_53 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  L0Memory_54 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  L0Memory_55 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  L0Memory_56 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  L0Memory_57 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  L0Memory_58 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  L0Memory_59 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  L0Memory_60 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  L0Memory_61 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  L0Memory_62 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  L0Memory_63 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  L0Memory_64 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  L0Memory_65 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  L0Memory_66 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  L0Memory_67 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  L0Memory_68 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  L0Memory_69 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  L0Memory_70 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  L0Memory_71 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  L0Memory_72 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  L0Memory_73 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  L0Memory_74 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  L0Memory_75 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  L0Memory_76 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  L0Memory_77 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  L0Memory_78 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  L0Memory_79 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  L0Memory_80 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  L0Memory_81 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  L0Memory_82 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  L0Memory_83 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  L0Memory_84 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  L0Memory_85 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  L0Memory_86 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  L0Memory_87 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  L0Memory_88 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  L0Memory_89 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  L0Memory_90 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  L0Memory_91 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  L0Memory_92 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  L0Memory_93 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  L0Memory_94 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  L0Memory_95 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  L0Memory_96 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  L0Memory_97 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  L0Memory_98 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  L0Memory_99 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  state = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  mux2out_reg = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  mux3out_reg = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  count = _RAND_104[9:0];
  _RAND_105 = {1{`RANDOM}};
  GRU_out_width = _RAND_105[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PE_22(
  input         clock,
  input         reset,
  input  [15:0] io_FromAbovePE,
  input  [15:0] io_FromLeftPE,
  input  [15:0] io_FromL1,
  input  [11:0] io_control_signal_mask,
  output [15:0] io_ToRightPE,
  output [15:0] io_ToBelowPE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] FP16MAC_io_a; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_b; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_c; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_out; // @[PEArray.scala 72:23]
  reg [5:0] L0Index; // @[PEArray.scala 39:24]
  reg [15:0] L0Memory_0; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_1; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_2; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_3; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_4; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_5; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_6; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_7; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_8; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_9; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_10; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_11; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_12; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_13; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_14; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_15; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_16; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_17; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_18; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_19; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_20; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_21; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_22; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_23; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_24; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_25; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_26; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_27; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_28; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_29; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_30; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_31; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_32; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_33; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_34; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_35; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_36; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_37; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_38; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_39; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_40; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_41; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_42; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_43; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_44; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_45; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_46; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_47; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_48; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_49; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_50; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_51; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_52; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_53; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_54; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_55; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_56; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_57; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_58; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_59; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_60; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_61; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_62; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_63; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_64; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_65; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_66; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_67; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_68; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_69; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_70; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_71; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_72; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_73; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_74; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_75; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_76; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_77; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_78; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_79; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_80; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_81; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_82; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_83; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_84; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_85; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_86; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_87; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_88; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_89; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_90; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_91; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_92; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_93; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_94; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_95; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_96; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_97; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_98; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_99; // @[PEArray.scala 40:21]
  reg [2:0] state; // @[PEArray.scala 100:22]
  wire  _T_3 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_12 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_16 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_22 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_31 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_41 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_342 = _T_41 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 231:12 PEArray.scala 32:8]
  wire  _GEN_349 = _T_31 ? 1'h0 : _GEN_342; // @[Conditional.scala 39:67 PEArray.scala 208:12]
  wire  _GEN_459 = _T_22 | _GEN_349; // @[Conditional.scala 39:67 PEArray.scala 32:8]
  wire  _GEN_463 = _T_16 ? 1'h0 : _GEN_459; // @[Conditional.scala 39:67]
  wire  _GEN_572 = _T_12 | _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 149:12]
  wire  sel1 = _T_3 | _GEN_572; // @[Conditional.scala 40:58 PEArray.scala 108:12]
  wire [15:0] MAC_out = FP16MAC_io_out; // @[PEArray.scala 47:21 PEArray.scala 85:11]
  wire  _GEN_465 = _T_16 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 177:12]
  wire  _GEN_580 = _T_12 | _GEN_465; // @[Conditional.scala 39:67 PEArray.scala 34:8]
  wire  sel3 = _T_3 | _GEN_580; // @[Conditional.scala 40:58 PEArray.scala 110:12]
  wire [1:0] _GEN_344 = _T_41 ? 2'h2 : 2'h0; // @[Conditional.scala 39:67 PEArray.scala 233:12 PEArray.scala 35:8]
  wire [1:0] _GEN_351 = _T_31 ? 2'h2 : _GEN_344; // @[Conditional.scala 39:67 PEArray.scala 210:12]
  wire [1:0] _GEN_461 = _T_22 ? 2'h0 : _GEN_351; // @[Conditional.scala 39:67 PEArray.scala 35:8]
  wire [1:0] _GEN_466 = _T_16 ? 2'h0 : _GEN_461; // @[Conditional.scala 39:67 PEArray.scala 178:12]
  wire [1:0] _GEN_574 = _T_12 ? 2'h1 : _GEN_466; // @[Conditional.scala 39:67]
  wire [1:0] sel4 = _T_3 ? 2'h0 : _GEN_574; // @[Conditional.scala 40:58 PEArray.scala 111:12]
  wire [15:0] _GEN_3 = sel4 == 2'h2 ? io_FromL1 : 16'h0; // @[PEArray.scala 65:28 PEArray.scala 66:15 PEArray.scala 69:15]
  wire [15:0] _GEN_4 = sel4 == 2'h1 ? io_FromAbovePE : _GEN_3; // @[PEArray.scala 62:28 PEArray.scala 63:15]
  wire [15:0] mux4out = sel4 == 2'h0 ? 16'h0 : _GEN_4; // @[PEArray.scala 59:22 PEArray.scala 60:13]
  wire [15:0] _GEN_7 = 6'h1 == L0Index ? L0Memory_1 : L0Memory_0; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_8 = 6'h2 == L0Index ? L0Memory_2 : _GEN_7; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_9 = 6'h3 == L0Index ? L0Memory_3 : _GEN_8; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_10 = 6'h4 == L0Index ? L0Memory_4 : _GEN_9; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_11 = 6'h5 == L0Index ? L0Memory_5 : _GEN_10; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_12 = 6'h6 == L0Index ? L0Memory_6 : _GEN_11; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_13 = 6'h7 == L0Index ? L0Memory_7 : _GEN_12; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_14 = 6'h8 == L0Index ? L0Memory_8 : _GEN_13; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_15 = 6'h9 == L0Index ? L0Memory_9 : _GEN_14; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_16 = 6'ha == L0Index ? L0Memory_10 : _GEN_15; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_17 = 6'hb == L0Index ? L0Memory_11 : _GEN_16; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_18 = 6'hc == L0Index ? L0Memory_12 : _GEN_17; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_19 = 6'hd == L0Index ? L0Memory_13 : _GEN_18; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_20 = 6'he == L0Index ? L0Memory_14 : _GEN_19; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_21 = 6'hf == L0Index ? L0Memory_15 : _GEN_20; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_22 = 6'h10 == L0Index ? L0Memory_16 : _GEN_21; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_23 = 6'h11 == L0Index ? L0Memory_17 : _GEN_22; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_24 = 6'h12 == L0Index ? L0Memory_18 : _GEN_23; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_25 = 6'h13 == L0Index ? L0Memory_19 : _GEN_24; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_26 = 6'h14 == L0Index ? L0Memory_20 : _GEN_25; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_27 = 6'h15 == L0Index ? L0Memory_21 : _GEN_26; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_28 = 6'h16 == L0Index ? L0Memory_22 : _GEN_27; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_29 = 6'h17 == L0Index ? L0Memory_23 : _GEN_28; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_30 = 6'h18 == L0Index ? L0Memory_24 : _GEN_29; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_31 = 6'h19 == L0Index ? L0Memory_25 : _GEN_30; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_32 = 6'h1a == L0Index ? L0Memory_26 : _GEN_31; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_33 = 6'h1b == L0Index ? L0Memory_27 : _GEN_32; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_34 = 6'h1c == L0Index ? L0Memory_28 : _GEN_33; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_35 = 6'h1d == L0Index ? L0Memory_29 : _GEN_34; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_36 = 6'h1e == L0Index ? L0Memory_30 : _GEN_35; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_37 = 6'h1f == L0Index ? L0Memory_31 : _GEN_36; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_38 = 6'h20 == L0Index ? L0Memory_32 : _GEN_37; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_39 = 6'h21 == L0Index ? L0Memory_33 : _GEN_38; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_40 = 6'h22 == L0Index ? L0Memory_34 : _GEN_39; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_41 = 6'h23 == L0Index ? L0Memory_35 : _GEN_40; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_42 = 6'h24 == L0Index ? L0Memory_36 : _GEN_41; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_43 = 6'h25 == L0Index ? L0Memory_37 : _GEN_42; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_44 = 6'h26 == L0Index ? L0Memory_38 : _GEN_43; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_45 = 6'h27 == L0Index ? L0Memory_39 : _GEN_44; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_46 = 6'h28 == L0Index ? L0Memory_40 : _GEN_45; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_47 = 6'h29 == L0Index ? L0Memory_41 : _GEN_46; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_48 = 6'h2a == L0Index ? L0Memory_42 : _GEN_47; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_49 = 6'h2b == L0Index ? L0Memory_43 : _GEN_48; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_50 = 6'h2c == L0Index ? L0Memory_44 : _GEN_49; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_51 = 6'h2d == L0Index ? L0Memory_45 : _GEN_50; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_52 = 6'h2e == L0Index ? L0Memory_46 : _GEN_51; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_53 = 6'h2f == L0Index ? L0Memory_47 : _GEN_52; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_54 = 6'h30 == L0Index ? L0Memory_48 : _GEN_53; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_55 = 6'h31 == L0Index ? L0Memory_49 : _GEN_54; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_56 = 6'h32 == L0Index ? L0Memory_50 : _GEN_55; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_57 = 6'h33 == L0Index ? L0Memory_51 : _GEN_56; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_58 = 6'h34 == L0Index ? L0Memory_52 : _GEN_57; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_59 = 6'h35 == L0Index ? L0Memory_53 : _GEN_58; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_60 = 6'h36 == L0Index ? L0Memory_54 : _GEN_59; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_61 = 6'h37 == L0Index ? L0Memory_55 : _GEN_60; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_62 = 6'h38 == L0Index ? L0Memory_56 : _GEN_61; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_63 = 6'h39 == L0Index ? L0Memory_57 : _GEN_62; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_64 = 6'h3a == L0Index ? L0Memory_58 : _GEN_63; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_65 = 6'h3b == L0Index ? L0Memory_59 : _GEN_64; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_66 = 6'h3c == L0Index ? L0Memory_60 : _GEN_65; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_67 = 6'h3d == L0Index ? L0Memory_61 : _GEN_66; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_68 = 6'h3e == L0Index ? L0Memory_62 : _GEN_67; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_69 = 6'h3f == L0Index ? L0Memory_63 : _GEN_68; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [6:0] _GEN_793 = {{1'd0}, L0Index}; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_70 = 7'h40 == _GEN_793 ? L0Memory_64 : _GEN_69; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_71 = 7'h41 == _GEN_793 ? L0Memory_65 : _GEN_70; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_72 = 7'h42 == _GEN_793 ? L0Memory_66 : _GEN_71; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_73 = 7'h43 == _GEN_793 ? L0Memory_67 : _GEN_72; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_74 = 7'h44 == _GEN_793 ? L0Memory_68 : _GEN_73; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_75 = 7'h45 == _GEN_793 ? L0Memory_69 : _GEN_74; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_76 = 7'h46 == _GEN_793 ? L0Memory_70 : _GEN_75; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_77 = 7'h47 == _GEN_793 ? L0Memory_71 : _GEN_76; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_78 = 7'h48 == _GEN_793 ? L0Memory_72 : _GEN_77; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_79 = 7'h49 == _GEN_793 ? L0Memory_73 : _GEN_78; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_80 = 7'h4a == _GEN_793 ? L0Memory_74 : _GEN_79; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_81 = 7'h4b == _GEN_793 ? L0Memory_75 : _GEN_80; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_82 = 7'h4c == _GEN_793 ? L0Memory_76 : _GEN_81; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_83 = 7'h4d == _GEN_793 ? L0Memory_77 : _GEN_82; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_84 = 7'h4e == _GEN_793 ? L0Memory_78 : _GEN_83; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_85 = 7'h4f == _GEN_793 ? L0Memory_79 : _GEN_84; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_86 = 7'h50 == _GEN_793 ? L0Memory_80 : _GEN_85; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_87 = 7'h51 == _GEN_793 ? L0Memory_81 : _GEN_86; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_88 = 7'h52 == _GEN_793 ? L0Memory_82 : _GEN_87; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_89 = 7'h53 == _GEN_793 ? L0Memory_83 : _GEN_88; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_90 = 7'h54 == _GEN_793 ? L0Memory_84 : _GEN_89; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_91 = 7'h55 == _GEN_793 ? L0Memory_85 : _GEN_90; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_92 = 7'h56 == _GEN_793 ? L0Memory_86 : _GEN_91; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_93 = 7'h57 == _GEN_793 ? L0Memory_87 : _GEN_92; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_94 = 7'h58 == _GEN_793 ? L0Memory_88 : _GEN_93; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_95 = 7'h59 == _GEN_793 ? L0Memory_89 : _GEN_94; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_96 = 7'h5a == _GEN_793 ? L0Memory_90 : _GEN_95; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_97 = 7'h5b == _GEN_793 ? L0Memory_91 : _GEN_96; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_98 = 7'h5c == _GEN_793 ? L0Memory_92 : _GEN_97; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_99 = 7'h5d == _GEN_793 ? L0Memory_93 : _GEN_98; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_100 = 7'h5e == _GEN_793 ? L0Memory_94 : _GEN_99; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_101 = 7'h5f == _GEN_793 ? L0Memory_95 : _GEN_100; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_102 = 7'h60 == _GEN_793 ? L0Memory_96 : _GEN_101; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_103 = 7'h61 == _GEN_793 ? L0Memory_97 : _GEN_102; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_104 = 7'h62 == _GEN_793 ? L0Memory_98 : _GEN_103; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_105 = 7'h63 == _GEN_793 ? L0Memory_99 : _GEN_104; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire  _GEN_575 = _T_12 ? 1'h0 : _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 157:12]
  wire  sel5 = _T_3 ? 1'h0 : _GEN_575; // @[Conditional.scala 40:58 PEArray.scala 112:12]
  reg [15:0] mux2out_reg; // @[PEArray.scala 90:28]
  reg [15:0] mux3out_reg; // @[PEArray.scala 91:28]
  reg [9:0] count; // @[PEArray.scala 101:22]
  reg [5:0] GRU_out_width; // @[PEArray.scala 104:26]
  wire [7:0] _GEN_118 = io_control_signal_mask[4] ? 8'h0 : {{2'd0}, GRU_out_width}; // @[PEArray.scala 116:57 PEArray.scala 145:23 PEArray.scala 104:26]
  wire [9:0] _count_T_1 = count + 10'h1; // @[PEArray.scala 162:24]
  wire [9:0] _GEN_120 = count != 10'h33 ? _count_T_1 : count; // @[PEArray.scala 161:27 PEArray.scala 162:15 PEArray.scala 101:22]
  wire [9:0] _GEN_124 = count != 10'h188 ? _count_T_1 : count; // @[PEArray.scala 183:28 PEArray.scala 184:15 PEArray.scala 101:22]
  wire [9:0] _GEN_125 = count == 10'h188 ? 10'h0 : _GEN_124; // @[PEArray.scala 186:28 PEArray.scala 187:15]
  wire [2:0] _GEN_126 = count == 10'h188 ? 3'h0 : state; // @[PEArray.scala 186:28 PEArray.scala 188:15 PEArray.scala 100:22]
  wire [9:0] _GEN_127 = count != 10'h0 ? _count_T_1 : count; // @[PEArray.scala 192:32 PEArray.scala 193:15 PEArray.scala 101:22]
  wire  _T_24 = count == 10'h0; // @[PEArray.scala 195:18]
  wire [5:0] _GEN_128 = count == 10'h0 ? 6'h0 : L0Index; // @[PEArray.scala 195:26 PEArray.scala 196:17 PEArray.scala 39:24]
  wire [9:0] _T_27 = 10'h0 - 10'h1; // @[PEArray.scala 198:51]
  wire [15:0] _GEN_129 = 6'h0 == L0Index ? io_FromL1 : L0Memory_0; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_130 = 6'h1 == L0Index ? io_FromL1 : L0Memory_1; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_131 = 6'h2 == L0Index ? io_FromL1 : L0Memory_2; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_132 = 6'h3 == L0Index ? io_FromL1 : L0Memory_3; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_133 = 6'h4 == L0Index ? io_FromL1 : L0Memory_4; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_134 = 6'h5 == L0Index ? io_FromL1 : L0Memory_5; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_135 = 6'h6 == L0Index ? io_FromL1 : L0Memory_6; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_136 = 6'h7 == L0Index ? io_FromL1 : L0Memory_7; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_137 = 6'h8 == L0Index ? io_FromL1 : L0Memory_8; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_138 = 6'h9 == L0Index ? io_FromL1 : L0Memory_9; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_139 = 6'ha == L0Index ? io_FromL1 : L0Memory_10; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_140 = 6'hb == L0Index ? io_FromL1 : L0Memory_11; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_141 = 6'hc == L0Index ? io_FromL1 : L0Memory_12; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_142 = 6'hd == L0Index ? io_FromL1 : L0Memory_13; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_143 = 6'he == L0Index ? io_FromL1 : L0Memory_14; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_144 = 6'hf == L0Index ? io_FromL1 : L0Memory_15; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_145 = 6'h10 == L0Index ? io_FromL1 : L0Memory_16; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_146 = 6'h11 == L0Index ? io_FromL1 : L0Memory_17; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_147 = 6'h12 == L0Index ? io_FromL1 : L0Memory_18; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_148 = 6'h13 == L0Index ? io_FromL1 : L0Memory_19; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_149 = 6'h14 == L0Index ? io_FromL1 : L0Memory_20; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_150 = 6'h15 == L0Index ? io_FromL1 : L0Memory_21; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_151 = 6'h16 == L0Index ? io_FromL1 : L0Memory_22; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_152 = 6'h17 == L0Index ? io_FromL1 : L0Memory_23; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_153 = 6'h18 == L0Index ? io_FromL1 : L0Memory_24; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_154 = 6'h19 == L0Index ? io_FromL1 : L0Memory_25; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_155 = 6'h1a == L0Index ? io_FromL1 : L0Memory_26; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_156 = 6'h1b == L0Index ? io_FromL1 : L0Memory_27; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_157 = 6'h1c == L0Index ? io_FromL1 : L0Memory_28; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_158 = 6'h1d == L0Index ? io_FromL1 : L0Memory_29; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_159 = 6'h1e == L0Index ? io_FromL1 : L0Memory_30; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_160 = 6'h1f == L0Index ? io_FromL1 : L0Memory_31; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_161 = 6'h20 == L0Index ? io_FromL1 : L0Memory_32; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_162 = 6'h21 == L0Index ? io_FromL1 : L0Memory_33; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_163 = 6'h22 == L0Index ? io_FromL1 : L0Memory_34; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_164 = 6'h23 == L0Index ? io_FromL1 : L0Memory_35; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_165 = 6'h24 == L0Index ? io_FromL1 : L0Memory_36; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_166 = 6'h25 == L0Index ? io_FromL1 : L0Memory_37; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_167 = 6'h26 == L0Index ? io_FromL1 : L0Memory_38; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_168 = 6'h27 == L0Index ? io_FromL1 : L0Memory_39; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_169 = 6'h28 == L0Index ? io_FromL1 : L0Memory_40; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_170 = 6'h29 == L0Index ? io_FromL1 : L0Memory_41; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_171 = 6'h2a == L0Index ? io_FromL1 : L0Memory_42; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_172 = 6'h2b == L0Index ? io_FromL1 : L0Memory_43; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_173 = 6'h2c == L0Index ? io_FromL1 : L0Memory_44; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_174 = 6'h2d == L0Index ? io_FromL1 : L0Memory_45; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_175 = 6'h2e == L0Index ? io_FromL1 : L0Memory_46; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_176 = 6'h2f == L0Index ? io_FromL1 : L0Memory_47; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_177 = 6'h30 == L0Index ? io_FromL1 : L0Memory_48; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_178 = 6'h31 == L0Index ? io_FromL1 : L0Memory_49; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_179 = 6'h32 == L0Index ? io_FromL1 : L0Memory_50; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_180 = 6'h33 == L0Index ? io_FromL1 : L0Memory_51; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_181 = 6'h34 == L0Index ? io_FromL1 : L0Memory_52; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_182 = 6'h35 == L0Index ? io_FromL1 : L0Memory_53; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_183 = 6'h36 == L0Index ? io_FromL1 : L0Memory_54; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_184 = 6'h37 == L0Index ? io_FromL1 : L0Memory_55; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_185 = 6'h38 == L0Index ? io_FromL1 : L0Memory_56; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_186 = 6'h39 == L0Index ? io_FromL1 : L0Memory_57; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_187 = 6'h3a == L0Index ? io_FromL1 : L0Memory_58; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_188 = 6'h3b == L0Index ? io_FromL1 : L0Memory_59; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_189 = 6'h3c == L0Index ? io_FromL1 : L0Memory_60; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_190 = 6'h3d == L0Index ? io_FromL1 : L0Memory_61; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_191 = 6'h3e == L0Index ? io_FromL1 : L0Memory_62; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_192 = 6'h3f == L0Index ? io_FromL1 : L0Memory_63; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_193 = 7'h40 == _GEN_793 ? io_FromL1 : L0Memory_64; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_194 = 7'h41 == _GEN_793 ? io_FromL1 : L0Memory_65; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_195 = 7'h42 == _GEN_793 ? io_FromL1 : L0Memory_66; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_196 = 7'h43 == _GEN_793 ? io_FromL1 : L0Memory_67; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_197 = 7'h44 == _GEN_793 ? io_FromL1 : L0Memory_68; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_198 = 7'h45 == _GEN_793 ? io_FromL1 : L0Memory_69; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_199 = 7'h46 == _GEN_793 ? io_FromL1 : L0Memory_70; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_200 = 7'h47 == _GEN_793 ? io_FromL1 : L0Memory_71; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_201 = 7'h48 == _GEN_793 ? io_FromL1 : L0Memory_72; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_202 = 7'h49 == _GEN_793 ? io_FromL1 : L0Memory_73; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_203 = 7'h4a == _GEN_793 ? io_FromL1 : L0Memory_74; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_204 = 7'h4b == _GEN_793 ? io_FromL1 : L0Memory_75; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_205 = 7'h4c == _GEN_793 ? io_FromL1 : L0Memory_76; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_206 = 7'h4d == _GEN_793 ? io_FromL1 : L0Memory_77; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_207 = 7'h4e == _GEN_793 ? io_FromL1 : L0Memory_78; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_208 = 7'h4f == _GEN_793 ? io_FromL1 : L0Memory_79; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_209 = 7'h50 == _GEN_793 ? io_FromL1 : L0Memory_80; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_210 = 7'h51 == _GEN_793 ? io_FromL1 : L0Memory_81; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_211 = 7'h52 == _GEN_793 ? io_FromL1 : L0Memory_82; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_212 = 7'h53 == _GEN_793 ? io_FromL1 : L0Memory_83; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_213 = 7'h54 == _GEN_793 ? io_FromL1 : L0Memory_84; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_214 = 7'h55 == _GEN_793 ? io_FromL1 : L0Memory_85; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_215 = 7'h56 == _GEN_793 ? io_FromL1 : L0Memory_86; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_216 = 7'h57 == _GEN_793 ? io_FromL1 : L0Memory_87; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_217 = 7'h58 == _GEN_793 ? io_FromL1 : L0Memory_88; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_218 = 7'h59 == _GEN_793 ? io_FromL1 : L0Memory_89; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_219 = 7'h5a == _GEN_793 ? io_FromL1 : L0Memory_90; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_220 = 7'h5b == _GEN_793 ? io_FromL1 : L0Memory_91; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_221 = 7'h5c == _GEN_793 ? io_FromL1 : L0Memory_92; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_222 = 7'h5d == _GEN_793 ? io_FromL1 : L0Memory_93; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_223 = 7'h5e == _GEN_793 ? io_FromL1 : L0Memory_94; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_224 = 7'h5f == _GEN_793 ? io_FromL1 : L0Memory_95; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_225 = 7'h60 == _GEN_793 ? io_FromL1 : L0Memory_96; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_226 = 7'h61 == _GEN_793 ? io_FromL1 : L0Memory_97; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_227 = 7'h62 == _GEN_793 ? io_FromL1 : L0Memory_98; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_228 = 7'h63 == _GEN_793 ? io_FromL1 : L0Memory_99; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [5:0] _L0Index_T_2 = L0Index + 6'h1; // @[PEArray.scala 200:28]
  wire [15:0] _GEN_229 = count >= 10'h1 & count <= _T_27 ? _GEN_129 : L0Memory_0; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_230 = count >= 10'h1 & count <= _T_27 ? _GEN_130 : L0Memory_1; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_231 = count >= 10'h1 & count <= _T_27 ? _GEN_131 : L0Memory_2; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_232 = count >= 10'h1 & count <= _T_27 ? _GEN_132 : L0Memory_3; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_233 = count >= 10'h1 & count <= _T_27 ? _GEN_133 : L0Memory_4; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_234 = count >= 10'h1 & count <= _T_27 ? _GEN_134 : L0Memory_5; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_235 = count >= 10'h1 & count <= _T_27 ? _GEN_135 : L0Memory_6; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_236 = count >= 10'h1 & count <= _T_27 ? _GEN_136 : L0Memory_7; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_237 = count >= 10'h1 & count <= _T_27 ? _GEN_137 : L0Memory_8; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_238 = count >= 10'h1 & count <= _T_27 ? _GEN_138 : L0Memory_9; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_239 = count >= 10'h1 & count <= _T_27 ? _GEN_139 : L0Memory_10; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_240 = count >= 10'h1 & count <= _T_27 ? _GEN_140 : L0Memory_11; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_241 = count >= 10'h1 & count <= _T_27 ? _GEN_141 : L0Memory_12; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_242 = count >= 10'h1 & count <= _T_27 ? _GEN_142 : L0Memory_13; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_243 = count >= 10'h1 & count <= _T_27 ? _GEN_143 : L0Memory_14; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_244 = count >= 10'h1 & count <= _T_27 ? _GEN_144 : L0Memory_15; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_245 = count >= 10'h1 & count <= _T_27 ? _GEN_145 : L0Memory_16; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_246 = count >= 10'h1 & count <= _T_27 ? _GEN_146 : L0Memory_17; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_247 = count >= 10'h1 & count <= _T_27 ? _GEN_147 : L0Memory_18; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_248 = count >= 10'h1 & count <= _T_27 ? _GEN_148 : L0Memory_19; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_249 = count >= 10'h1 & count <= _T_27 ? _GEN_149 : L0Memory_20; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_250 = count >= 10'h1 & count <= _T_27 ? _GEN_150 : L0Memory_21; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_251 = count >= 10'h1 & count <= _T_27 ? _GEN_151 : L0Memory_22; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_252 = count >= 10'h1 & count <= _T_27 ? _GEN_152 : L0Memory_23; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_253 = count >= 10'h1 & count <= _T_27 ? _GEN_153 : L0Memory_24; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_254 = count >= 10'h1 & count <= _T_27 ? _GEN_154 : L0Memory_25; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_255 = count >= 10'h1 & count <= _T_27 ? _GEN_155 : L0Memory_26; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_256 = count >= 10'h1 & count <= _T_27 ? _GEN_156 : L0Memory_27; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_257 = count >= 10'h1 & count <= _T_27 ? _GEN_157 : L0Memory_28; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_258 = count >= 10'h1 & count <= _T_27 ? _GEN_158 : L0Memory_29; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_259 = count >= 10'h1 & count <= _T_27 ? _GEN_159 : L0Memory_30; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_260 = count >= 10'h1 & count <= _T_27 ? _GEN_160 : L0Memory_31; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_261 = count >= 10'h1 & count <= _T_27 ? _GEN_161 : L0Memory_32; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_262 = count >= 10'h1 & count <= _T_27 ? _GEN_162 : L0Memory_33; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_263 = count >= 10'h1 & count <= _T_27 ? _GEN_163 : L0Memory_34; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_264 = count >= 10'h1 & count <= _T_27 ? _GEN_164 : L0Memory_35; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_265 = count >= 10'h1 & count <= _T_27 ? _GEN_165 : L0Memory_36; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_266 = count >= 10'h1 & count <= _T_27 ? _GEN_166 : L0Memory_37; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_267 = count >= 10'h1 & count <= _T_27 ? _GEN_167 : L0Memory_38; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_268 = count >= 10'h1 & count <= _T_27 ? _GEN_168 : L0Memory_39; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_269 = count >= 10'h1 & count <= _T_27 ? _GEN_169 : L0Memory_40; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_270 = count >= 10'h1 & count <= _T_27 ? _GEN_170 : L0Memory_41; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_271 = count >= 10'h1 & count <= _T_27 ? _GEN_171 : L0Memory_42; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_272 = count >= 10'h1 & count <= _T_27 ? _GEN_172 : L0Memory_43; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_273 = count >= 10'h1 & count <= _T_27 ? _GEN_173 : L0Memory_44; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_274 = count >= 10'h1 & count <= _T_27 ? _GEN_174 : L0Memory_45; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_275 = count >= 10'h1 & count <= _T_27 ? _GEN_175 : L0Memory_46; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_276 = count >= 10'h1 & count <= _T_27 ? _GEN_176 : L0Memory_47; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_277 = count >= 10'h1 & count <= _T_27 ? _GEN_177 : L0Memory_48; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_278 = count >= 10'h1 & count <= _T_27 ? _GEN_178 : L0Memory_49; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_279 = count >= 10'h1 & count <= _T_27 ? _GEN_179 : L0Memory_50; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_280 = count >= 10'h1 & count <= _T_27 ? _GEN_180 : L0Memory_51; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_281 = count >= 10'h1 & count <= _T_27 ? _GEN_181 : L0Memory_52; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_282 = count >= 10'h1 & count <= _T_27 ? _GEN_182 : L0Memory_53; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_283 = count >= 10'h1 & count <= _T_27 ? _GEN_183 : L0Memory_54; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_284 = count >= 10'h1 & count <= _T_27 ? _GEN_184 : L0Memory_55; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_285 = count >= 10'h1 & count <= _T_27 ? _GEN_185 : L0Memory_56; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_286 = count >= 10'h1 & count <= _T_27 ? _GEN_186 : L0Memory_57; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_287 = count >= 10'h1 & count <= _T_27 ? _GEN_187 : L0Memory_58; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_288 = count >= 10'h1 & count <= _T_27 ? _GEN_188 : L0Memory_59; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_289 = count >= 10'h1 & count <= _T_27 ? _GEN_189 : L0Memory_60; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_290 = count >= 10'h1 & count <= _T_27 ? _GEN_190 : L0Memory_61; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_291 = count >= 10'h1 & count <= _T_27 ? _GEN_191 : L0Memory_62; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_292 = count >= 10'h1 & count <= _T_27 ? _GEN_192 : L0Memory_63; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_293 = count >= 10'h1 & count <= _T_27 ? _GEN_193 : L0Memory_64; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_294 = count >= 10'h1 & count <= _T_27 ? _GEN_194 : L0Memory_65; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_295 = count >= 10'h1 & count <= _T_27 ? _GEN_195 : L0Memory_66; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_296 = count >= 10'h1 & count <= _T_27 ? _GEN_196 : L0Memory_67; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_297 = count >= 10'h1 & count <= _T_27 ? _GEN_197 : L0Memory_68; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_298 = count >= 10'h1 & count <= _T_27 ? _GEN_198 : L0Memory_69; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_299 = count >= 10'h1 & count <= _T_27 ? _GEN_199 : L0Memory_70; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_300 = count >= 10'h1 & count <= _T_27 ? _GEN_200 : L0Memory_71; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_301 = count >= 10'h1 & count <= _T_27 ? _GEN_201 : L0Memory_72; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_302 = count >= 10'h1 & count <= _T_27 ? _GEN_202 : L0Memory_73; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_303 = count >= 10'h1 & count <= _T_27 ? _GEN_203 : L0Memory_74; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_304 = count >= 10'h1 & count <= _T_27 ? _GEN_204 : L0Memory_75; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_305 = count >= 10'h1 & count <= _T_27 ? _GEN_205 : L0Memory_76; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_306 = count >= 10'h1 & count <= _T_27 ? _GEN_206 : L0Memory_77; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_307 = count >= 10'h1 & count <= _T_27 ? _GEN_207 : L0Memory_78; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_308 = count >= 10'h1 & count <= _T_27 ? _GEN_208 : L0Memory_79; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_309 = count >= 10'h1 & count <= _T_27 ? _GEN_209 : L0Memory_80; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_310 = count >= 10'h1 & count <= _T_27 ? _GEN_210 : L0Memory_81; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_311 = count >= 10'h1 & count <= _T_27 ? _GEN_211 : L0Memory_82; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_312 = count >= 10'h1 & count <= _T_27 ? _GEN_212 : L0Memory_83; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_313 = count >= 10'h1 & count <= _T_27 ? _GEN_213 : L0Memory_84; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_314 = count >= 10'h1 & count <= _T_27 ? _GEN_214 : L0Memory_85; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_315 = count >= 10'h1 & count <= _T_27 ? _GEN_215 : L0Memory_86; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_316 = count >= 10'h1 & count <= _T_27 ? _GEN_216 : L0Memory_87; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_317 = count >= 10'h1 & count <= _T_27 ? _GEN_217 : L0Memory_88; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_318 = count >= 10'h1 & count <= _T_27 ? _GEN_218 : L0Memory_89; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_319 = count >= 10'h1 & count <= _T_27 ? _GEN_219 : L0Memory_90; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_320 = count >= 10'h1 & count <= _T_27 ? _GEN_220 : L0Memory_91; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_321 = count >= 10'h1 & count <= _T_27 ? _GEN_221 : L0Memory_92; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_322 = count >= 10'h1 & count <= _T_27 ? _GEN_222 : L0Memory_93; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_323 = count >= 10'h1 & count <= _T_27 ? _GEN_223 : L0Memory_94; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_324 = count >= 10'h1 & count <= _T_27 ? _GEN_224 : L0Memory_95; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_325 = count >= 10'h1 & count <= _T_27 ? _GEN_225 : L0Memory_96; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_326 = count >= 10'h1 & count <= _T_27 ? _GEN_226 : L0Memory_97; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_327 = count >= 10'h1 & count <= _T_27 ? _GEN_227 : L0Memory_98; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_328 = count >= 10'h1 & count <= _T_27 ? _GEN_228 : L0Memory_99; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [5:0] _GEN_329 = count >= 10'h1 & count <= _T_27 ? _L0Index_T_2 : _GEN_128; // @[PEArray.scala 198:59 PEArray.scala 200:17]
  wire [9:0] _GEN_330 = _T_24 ? 10'h0 : _GEN_127; // @[PEArray.scala 202:32 PEArray.scala 203:15]
  wire [2:0] _GEN_331 = _T_24 ? 3'h0 : state; // @[PEArray.scala 202:32 PEArray.scala 204:15 PEArray.scala 100:22]
  wire [9:0] _GEN_865 = {{4'd0}, GRU_out_width}; // @[PEArray.scala 220:19]
  wire [9:0] _GEN_0 = count % _GEN_865; // @[PEArray.scala 220:19]
  wire [5:0] _T_36 = _GEN_0[5:0]; // @[PEArray.scala 220:19]
  wire [5:0] _T_38 = GRU_out_width - 6'h1; // @[PEArray.scala 220:55]
  wire [5:0] _GEN_334 = _T_36 == _T_38 ? _L0Index_T_2 : 6'h0; // @[PEArray.scala 220:62 PEArray.scala 221:17 PEArray.scala 214:15]
  wire [5:0] _GEN_346 = _T_41 ? _GEN_334 : L0Index; // @[Conditional.scala 39:67 PEArray.scala 39:24]
  wire [9:0] _GEN_347 = _T_41 ? _GEN_330 : count; // @[Conditional.scala 39:67 PEArray.scala 101:22]
  wire [2:0] _GEN_348 = _T_41 ? _GEN_331 : state; // @[Conditional.scala 39:67 PEArray.scala 100:22]
  wire [5:0] _GEN_353 = _T_31 ? _GEN_334 : _GEN_346; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_354 = _T_31 ? _GEN_330 : _GEN_347; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_355 = _T_31 ? _GEN_331 : _GEN_348; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_356 = _T_22 ? _GEN_330 : _GEN_354; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_357 = _T_22 ? _GEN_329 : _GEN_353; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_458 = _T_22 ? _GEN_331 : _GEN_355; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_690 = _T_3 ? _GEN_118 : {{2'd0}, GRU_out_width}; // @[Conditional.scala 40:58 PEArray.scala 104:26]
  FP16MulAdder FP16MAC ( // @[PEArray.scala 72:23]
    .io_a(FP16MAC_io_a),
    .io_b(FP16MAC_io_b),
    .io_c(FP16MAC_io_c),
    .io_out(FP16MAC_io_out)
  );
  assign io_ToRightPE = mux3out_reg; // @[PEArray.scala 95:16]
  assign io_ToBelowPE = mux2out_reg; // @[PEArray.scala 94:16]
  assign FP16MAC_io_a = sel1 ? io_FromL1 : io_FromLeftPE; // @[PEArray.scala 50:14 PEArray.scala 50:23 PEArray.scala 51:24]
  assign FP16MAC_io_b = sel5 ? mux4out : _GEN_105; // @[PEArray.scala 77:13 PEArray.scala 78:18 PEArray.scala 81:18]
  assign FP16MAC_io_c = sel5 ? _GEN_105 : mux4out; // @[PEArray.scala 77:13 PEArray.scala 79:18 PEArray.scala 82:18]
  always @(posedge clock) begin
    if (reset) begin // @[PEArray.scala 39:24]
      L0Index <= 6'h0; // @[PEArray.scala 39:24]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h1; // @[PEArray.scala 159:15]
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        L0Index <= 6'ha; // @[PEArray.scala 181:15]
      end else begin
        L0Index <= _GEN_357;
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_0 <= _GEN_229;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_1 <= _GEN_230;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_2 <= _GEN_231;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_3 <= _GEN_232;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_4 <= _GEN_233;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_5 <= _GEN_234;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_6 <= _GEN_235;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_7 <= _GEN_236;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_8 <= _GEN_237;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_9 <= _GEN_238;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_10 <= _GEN_239;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_11 <= _GEN_240;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_12 <= _GEN_241;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_13 <= _GEN_242;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_14 <= _GEN_243;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_15 <= _GEN_244;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_16 <= _GEN_245;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_17 <= _GEN_246;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_18 <= _GEN_247;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_19 <= _GEN_248;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_20 <= _GEN_249;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_21 <= _GEN_250;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_22 <= _GEN_251;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_23 <= _GEN_252;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_24 <= _GEN_253;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_25 <= _GEN_254;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_26 <= _GEN_255;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_27 <= _GEN_256;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_28 <= _GEN_257;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_29 <= _GEN_258;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_30 <= _GEN_259;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_31 <= _GEN_260;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_32 <= _GEN_261;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_33 <= _GEN_262;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_34 <= _GEN_263;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_35 <= _GEN_264;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_36 <= _GEN_265;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_37 <= _GEN_266;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_38 <= _GEN_267;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_39 <= _GEN_268;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_40 <= _GEN_269;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_41 <= _GEN_270;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_42 <= _GEN_271;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_43 <= _GEN_272;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_44 <= _GEN_273;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_45 <= _GEN_274;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_46 <= _GEN_275;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_47 <= _GEN_276;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_48 <= _GEN_277;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_49 <= _GEN_278;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_50 <= _GEN_279;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_51 <= _GEN_280;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_52 <= _GEN_281;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_53 <= _GEN_282;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_54 <= _GEN_283;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_55 <= _GEN_284;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_56 <= _GEN_285;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_57 <= _GEN_286;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_58 <= _GEN_287;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_59 <= _GEN_288;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_60 <= _GEN_289;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_61 <= _GEN_290;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_62 <= _GEN_291;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_63 <= _GEN_292;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_64 <= _GEN_293;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_65 <= _GEN_294;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_66 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_67 <= _GEN_296;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_68 <= _GEN_297;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_69 <= _GEN_298;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_70 <= _GEN_299;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_71 <= _GEN_300;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_72 <= _GEN_301;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_73 <= _GEN_302;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_74 <= _GEN_303;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_75 <= _GEN_304;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_76 <= _GEN_305;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_77 <= _GEN_306;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_78 <= _GEN_307;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_79 <= _GEN_308;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_80 <= _GEN_309;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_81 <= _GEN_310;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_82 <= _GEN_311;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_83 <= _GEN_312;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_84 <= _GEN_313;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_85 <= _GEN_314;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_86 <= _GEN_315;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_87 <= _GEN_316;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_88 <= _GEN_317;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_89 <= _GEN_318;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_90 <= _GEN_319;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_91 <= _GEN_320;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_92 <= _GEN_321;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_93 <= _GEN_322;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_94 <= _GEN_323;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_95 <= _GEN_324;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_96 <= _GEN_325;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_97 <= _GEN_326;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_98 <= _GEN_327;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_99 <= _GEN_328;
          end
        end
      end
    end
    if (reset) begin // @[PEArray.scala 100:22]
      state <= 3'h0; // @[PEArray.scala 100:22]
    end else if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[4]) begin // @[PEArray.scala 116:57]
        state <= 3'h1;
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      if (count == 10'h33) begin // @[PEArray.scala 164:27]
        state <= 3'h0; // @[PEArray.scala 166:15]
      end
    end else if (_T_16) begin // @[Conditional.scala 39:67]
      state <= _GEN_126;
    end else begin
      state <= _GEN_458;
    end
    if (reset) begin // @[PEArray.scala 90:28]
      mux2out_reg <= 16'h0; // @[PEArray.scala 90:28]
    end else begin
      mux2out_reg <= MAC_out; // @[PEArray.scala 90:28]
    end
    if (reset) begin // @[PEArray.scala 91:28]
      mux3out_reg <= 16'h0; // @[PEArray.scala 91:28]
    end else if (sel3) begin // @[PEArray.scala 56:14]
      mux3out_reg <= MAC_out; // @[PEArray.scala 56:23]
    end else if (sel1) begin // @[PEArray.scala 50:14]
      mux3out_reg <= io_FromL1; // @[PEArray.scala 50:23]
    end else begin
      mux3out_reg <= io_FromLeftPE; // @[PEArray.scala 51:24]
    end
    if (reset) begin // @[PEArray.scala 101:22]
      count <= 10'h0; // @[PEArray.scala 101:22]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        if (count == 10'h33) begin // @[PEArray.scala 164:27]
          count <= 10'h0; // @[PEArray.scala 165:15]
        end else begin
          count <= _GEN_120;
        end
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        count <= _GEN_125;
      end else begin
        count <= _GEN_356;
      end
    end
    GRU_out_width <= _GEN_690[5:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  L0Index = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  L0Memory_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  L0Memory_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  L0Memory_2 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  L0Memory_3 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  L0Memory_4 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  L0Memory_5 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  L0Memory_6 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  L0Memory_7 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  L0Memory_8 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  L0Memory_9 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  L0Memory_10 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  L0Memory_11 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  L0Memory_12 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  L0Memory_13 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  L0Memory_14 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  L0Memory_15 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  L0Memory_16 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  L0Memory_17 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  L0Memory_18 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  L0Memory_19 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  L0Memory_20 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  L0Memory_21 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  L0Memory_22 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  L0Memory_23 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  L0Memory_24 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  L0Memory_25 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  L0Memory_26 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  L0Memory_27 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  L0Memory_28 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  L0Memory_29 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  L0Memory_30 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  L0Memory_31 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  L0Memory_32 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  L0Memory_33 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  L0Memory_34 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  L0Memory_35 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  L0Memory_36 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  L0Memory_37 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  L0Memory_38 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  L0Memory_39 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  L0Memory_40 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  L0Memory_41 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  L0Memory_42 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  L0Memory_43 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  L0Memory_44 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  L0Memory_45 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  L0Memory_46 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  L0Memory_47 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  L0Memory_48 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  L0Memory_49 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  L0Memory_50 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  L0Memory_51 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  L0Memory_52 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  L0Memory_53 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  L0Memory_54 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  L0Memory_55 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  L0Memory_56 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  L0Memory_57 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  L0Memory_58 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  L0Memory_59 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  L0Memory_60 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  L0Memory_61 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  L0Memory_62 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  L0Memory_63 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  L0Memory_64 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  L0Memory_65 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  L0Memory_66 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  L0Memory_67 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  L0Memory_68 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  L0Memory_69 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  L0Memory_70 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  L0Memory_71 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  L0Memory_72 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  L0Memory_73 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  L0Memory_74 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  L0Memory_75 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  L0Memory_76 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  L0Memory_77 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  L0Memory_78 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  L0Memory_79 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  L0Memory_80 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  L0Memory_81 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  L0Memory_82 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  L0Memory_83 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  L0Memory_84 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  L0Memory_85 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  L0Memory_86 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  L0Memory_87 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  L0Memory_88 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  L0Memory_89 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  L0Memory_90 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  L0Memory_91 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  L0Memory_92 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  L0Memory_93 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  L0Memory_94 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  L0Memory_95 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  L0Memory_96 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  L0Memory_97 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  L0Memory_98 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  L0Memory_99 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  state = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  mux2out_reg = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  mux3out_reg = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  count = _RAND_104[9:0];
  _RAND_105 = {1{`RANDOM}};
  GRU_out_width = _RAND_105[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PE_23(
  input         clock,
  input         reset,
  input  [15:0] io_FromAbovePE,
  input  [15:0] io_FromLeftPE,
  input  [15:0] io_FromL1,
  input  [2:0]  io_control_signal_control,
  input  [9:0]  io_control_signal_count,
  input  [5:0]  io_control_signal_L0index,
  input  [11:0] io_control_signal_mask,
  input  [7:0]  io_control_signal_gru_out_width,
  output [15:0] io_ToRightPE,
  output [15:0] io_ToBelowPE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] FP16MAC_io_a; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_b; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_c; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_out; // @[PEArray.scala 72:23]
  reg [5:0] L0Index; // @[PEArray.scala 39:24]
  reg [15:0] L0Memory_0; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_1; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_2; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_3; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_4; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_5; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_6; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_7; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_8; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_9; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_10; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_11; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_12; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_13; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_14; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_15; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_16; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_17; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_18; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_19; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_20; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_21; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_22; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_23; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_24; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_25; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_26; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_27; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_28; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_29; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_30; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_31; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_32; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_33; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_34; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_35; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_36; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_37; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_38; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_39; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_40; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_41; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_42; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_43; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_44; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_45; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_46; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_47; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_48; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_49; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_50; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_51; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_52; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_53; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_54; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_55; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_56; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_57; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_58; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_59; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_60; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_61; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_62; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_63; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_64; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_65; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_66; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_67; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_68; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_69; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_70; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_71; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_72; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_73; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_74; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_75; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_76; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_77; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_78; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_79; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_80; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_81; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_82; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_83; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_84; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_85; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_86; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_87; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_88; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_89; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_90; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_91; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_92; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_93; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_94; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_95; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_96; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_97; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_98; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_99; // @[PEArray.scala 40:21]
  reg [2:0] state; // @[PEArray.scala 100:22]
  wire  _T_3 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_12 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_16 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_22 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_31 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_41 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_342 = _T_41 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 231:12 PEArray.scala 32:8]
  wire  _GEN_349 = _T_31 ? 1'h0 : _GEN_342; // @[Conditional.scala 39:67 PEArray.scala 208:12]
  wire  _GEN_459 = _T_22 | _GEN_349; // @[Conditional.scala 39:67 PEArray.scala 32:8]
  wire  _GEN_463 = _T_16 ? 1'h0 : _GEN_459; // @[Conditional.scala 39:67]
  wire  _GEN_572 = _T_12 | _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 149:12]
  wire  sel1 = _T_3 | _GEN_572; // @[Conditional.scala 40:58 PEArray.scala 108:12]
  wire [15:0] MAC_out = FP16MAC_io_out; // @[PEArray.scala 47:21 PEArray.scala 85:11]
  wire  _GEN_465 = _T_16 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 177:12]
  wire  _GEN_580 = _T_12 | _GEN_465; // @[Conditional.scala 39:67 PEArray.scala 34:8]
  wire  sel3 = _T_3 | _GEN_580; // @[Conditional.scala 40:58 PEArray.scala 110:12]
  wire [1:0] _GEN_344 = _T_41 ? 2'h2 : 2'h0; // @[Conditional.scala 39:67 PEArray.scala 233:12 PEArray.scala 35:8]
  wire [1:0] _GEN_351 = _T_31 ? 2'h2 : _GEN_344; // @[Conditional.scala 39:67 PEArray.scala 210:12]
  wire [1:0] _GEN_461 = _T_22 ? 2'h0 : _GEN_351; // @[Conditional.scala 39:67 PEArray.scala 35:8]
  wire [1:0] _GEN_466 = _T_16 ? 2'h0 : _GEN_461; // @[Conditional.scala 39:67 PEArray.scala 178:12]
  wire [1:0] _GEN_574 = _T_12 ? 2'h1 : _GEN_466; // @[Conditional.scala 39:67]
  wire [1:0] sel4 = _T_3 ? 2'h0 : _GEN_574; // @[Conditional.scala 40:58 PEArray.scala 111:12]
  wire [15:0] _GEN_3 = sel4 == 2'h2 ? io_FromL1 : 16'h0; // @[PEArray.scala 65:28 PEArray.scala 66:15 PEArray.scala 69:15]
  wire [15:0] _GEN_4 = sel4 == 2'h1 ? io_FromAbovePE : _GEN_3; // @[PEArray.scala 62:28 PEArray.scala 63:15]
  wire [15:0] mux4out = sel4 == 2'h0 ? 16'h0 : _GEN_4; // @[PEArray.scala 59:22 PEArray.scala 60:13]
  wire [15:0] _GEN_7 = 6'h1 == L0Index ? L0Memory_1 : L0Memory_0; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_8 = 6'h2 == L0Index ? L0Memory_2 : _GEN_7; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_9 = 6'h3 == L0Index ? L0Memory_3 : _GEN_8; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_10 = 6'h4 == L0Index ? L0Memory_4 : _GEN_9; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_11 = 6'h5 == L0Index ? L0Memory_5 : _GEN_10; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_12 = 6'h6 == L0Index ? L0Memory_6 : _GEN_11; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_13 = 6'h7 == L0Index ? L0Memory_7 : _GEN_12; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_14 = 6'h8 == L0Index ? L0Memory_8 : _GEN_13; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_15 = 6'h9 == L0Index ? L0Memory_9 : _GEN_14; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_16 = 6'ha == L0Index ? L0Memory_10 : _GEN_15; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_17 = 6'hb == L0Index ? L0Memory_11 : _GEN_16; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_18 = 6'hc == L0Index ? L0Memory_12 : _GEN_17; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_19 = 6'hd == L0Index ? L0Memory_13 : _GEN_18; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_20 = 6'he == L0Index ? L0Memory_14 : _GEN_19; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_21 = 6'hf == L0Index ? L0Memory_15 : _GEN_20; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_22 = 6'h10 == L0Index ? L0Memory_16 : _GEN_21; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_23 = 6'h11 == L0Index ? L0Memory_17 : _GEN_22; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_24 = 6'h12 == L0Index ? L0Memory_18 : _GEN_23; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_25 = 6'h13 == L0Index ? L0Memory_19 : _GEN_24; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_26 = 6'h14 == L0Index ? L0Memory_20 : _GEN_25; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_27 = 6'h15 == L0Index ? L0Memory_21 : _GEN_26; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_28 = 6'h16 == L0Index ? L0Memory_22 : _GEN_27; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_29 = 6'h17 == L0Index ? L0Memory_23 : _GEN_28; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_30 = 6'h18 == L0Index ? L0Memory_24 : _GEN_29; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_31 = 6'h19 == L0Index ? L0Memory_25 : _GEN_30; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_32 = 6'h1a == L0Index ? L0Memory_26 : _GEN_31; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_33 = 6'h1b == L0Index ? L0Memory_27 : _GEN_32; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_34 = 6'h1c == L0Index ? L0Memory_28 : _GEN_33; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_35 = 6'h1d == L0Index ? L0Memory_29 : _GEN_34; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_36 = 6'h1e == L0Index ? L0Memory_30 : _GEN_35; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_37 = 6'h1f == L0Index ? L0Memory_31 : _GEN_36; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_38 = 6'h20 == L0Index ? L0Memory_32 : _GEN_37; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_39 = 6'h21 == L0Index ? L0Memory_33 : _GEN_38; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_40 = 6'h22 == L0Index ? L0Memory_34 : _GEN_39; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_41 = 6'h23 == L0Index ? L0Memory_35 : _GEN_40; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_42 = 6'h24 == L0Index ? L0Memory_36 : _GEN_41; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_43 = 6'h25 == L0Index ? L0Memory_37 : _GEN_42; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_44 = 6'h26 == L0Index ? L0Memory_38 : _GEN_43; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_45 = 6'h27 == L0Index ? L0Memory_39 : _GEN_44; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_46 = 6'h28 == L0Index ? L0Memory_40 : _GEN_45; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_47 = 6'h29 == L0Index ? L0Memory_41 : _GEN_46; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_48 = 6'h2a == L0Index ? L0Memory_42 : _GEN_47; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_49 = 6'h2b == L0Index ? L0Memory_43 : _GEN_48; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_50 = 6'h2c == L0Index ? L0Memory_44 : _GEN_49; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_51 = 6'h2d == L0Index ? L0Memory_45 : _GEN_50; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_52 = 6'h2e == L0Index ? L0Memory_46 : _GEN_51; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_53 = 6'h2f == L0Index ? L0Memory_47 : _GEN_52; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_54 = 6'h30 == L0Index ? L0Memory_48 : _GEN_53; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_55 = 6'h31 == L0Index ? L0Memory_49 : _GEN_54; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_56 = 6'h32 == L0Index ? L0Memory_50 : _GEN_55; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_57 = 6'h33 == L0Index ? L0Memory_51 : _GEN_56; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_58 = 6'h34 == L0Index ? L0Memory_52 : _GEN_57; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_59 = 6'h35 == L0Index ? L0Memory_53 : _GEN_58; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_60 = 6'h36 == L0Index ? L0Memory_54 : _GEN_59; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_61 = 6'h37 == L0Index ? L0Memory_55 : _GEN_60; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_62 = 6'h38 == L0Index ? L0Memory_56 : _GEN_61; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_63 = 6'h39 == L0Index ? L0Memory_57 : _GEN_62; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_64 = 6'h3a == L0Index ? L0Memory_58 : _GEN_63; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_65 = 6'h3b == L0Index ? L0Memory_59 : _GEN_64; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_66 = 6'h3c == L0Index ? L0Memory_60 : _GEN_65; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_67 = 6'h3d == L0Index ? L0Memory_61 : _GEN_66; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_68 = 6'h3e == L0Index ? L0Memory_62 : _GEN_67; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_69 = 6'h3f == L0Index ? L0Memory_63 : _GEN_68; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [6:0] _GEN_793 = {{1'd0}, L0Index}; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_70 = 7'h40 == _GEN_793 ? L0Memory_64 : _GEN_69; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_71 = 7'h41 == _GEN_793 ? L0Memory_65 : _GEN_70; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_72 = 7'h42 == _GEN_793 ? L0Memory_66 : _GEN_71; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_73 = 7'h43 == _GEN_793 ? L0Memory_67 : _GEN_72; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_74 = 7'h44 == _GEN_793 ? L0Memory_68 : _GEN_73; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_75 = 7'h45 == _GEN_793 ? L0Memory_69 : _GEN_74; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_76 = 7'h46 == _GEN_793 ? L0Memory_70 : _GEN_75; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_77 = 7'h47 == _GEN_793 ? L0Memory_71 : _GEN_76; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_78 = 7'h48 == _GEN_793 ? L0Memory_72 : _GEN_77; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_79 = 7'h49 == _GEN_793 ? L0Memory_73 : _GEN_78; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_80 = 7'h4a == _GEN_793 ? L0Memory_74 : _GEN_79; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_81 = 7'h4b == _GEN_793 ? L0Memory_75 : _GEN_80; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_82 = 7'h4c == _GEN_793 ? L0Memory_76 : _GEN_81; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_83 = 7'h4d == _GEN_793 ? L0Memory_77 : _GEN_82; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_84 = 7'h4e == _GEN_793 ? L0Memory_78 : _GEN_83; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_85 = 7'h4f == _GEN_793 ? L0Memory_79 : _GEN_84; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_86 = 7'h50 == _GEN_793 ? L0Memory_80 : _GEN_85; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_87 = 7'h51 == _GEN_793 ? L0Memory_81 : _GEN_86; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_88 = 7'h52 == _GEN_793 ? L0Memory_82 : _GEN_87; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_89 = 7'h53 == _GEN_793 ? L0Memory_83 : _GEN_88; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_90 = 7'h54 == _GEN_793 ? L0Memory_84 : _GEN_89; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_91 = 7'h55 == _GEN_793 ? L0Memory_85 : _GEN_90; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_92 = 7'h56 == _GEN_793 ? L0Memory_86 : _GEN_91; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_93 = 7'h57 == _GEN_793 ? L0Memory_87 : _GEN_92; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_94 = 7'h58 == _GEN_793 ? L0Memory_88 : _GEN_93; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_95 = 7'h59 == _GEN_793 ? L0Memory_89 : _GEN_94; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_96 = 7'h5a == _GEN_793 ? L0Memory_90 : _GEN_95; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_97 = 7'h5b == _GEN_793 ? L0Memory_91 : _GEN_96; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_98 = 7'h5c == _GEN_793 ? L0Memory_92 : _GEN_97; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_99 = 7'h5d == _GEN_793 ? L0Memory_93 : _GEN_98; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_100 = 7'h5e == _GEN_793 ? L0Memory_94 : _GEN_99; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_101 = 7'h5f == _GEN_793 ? L0Memory_95 : _GEN_100; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_102 = 7'h60 == _GEN_793 ? L0Memory_96 : _GEN_101; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_103 = 7'h61 == _GEN_793 ? L0Memory_97 : _GEN_102; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_104 = 7'h62 == _GEN_793 ? L0Memory_98 : _GEN_103; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_105 = 7'h63 == _GEN_793 ? L0Memory_99 : _GEN_104; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire  _GEN_575 = _T_12 ? 1'h0 : _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 157:12]
  wire  sel5 = _T_3 ? 1'h0 : _GEN_575; // @[Conditional.scala 40:58 PEArray.scala 112:12]
  reg [15:0] mux2out_reg; // @[PEArray.scala 90:28]
  reg [15:0] mux3out_reg; // @[PEArray.scala 91:28]
  reg [9:0] count; // @[PEArray.scala 101:22]
  reg [9:0] count_max; // @[PEArray.scala 102:22]
  reg [5:0] L0index_begin; // @[PEArray.scala 103:26]
  reg [5:0] GRU_out_width; // @[PEArray.scala 104:26]
  wire  _T_6 = 3'h0 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_7 = 3'h1 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_8 = 3'h2 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_9 = 3'h3 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_10 = 3'h4 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_11 = 3'h5 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_109 = _T_11 ? 3'h5 : state; // @[Conditional.scala 39:67 PEArray.scala 140:19 PEArray.scala 100:22]
  wire [2:0] _GEN_110 = _T_10 ? 3'h4 : _GEN_109; // @[Conditional.scala 39:67 PEArray.scala 136:19]
  wire [2:0] _GEN_111 = _T_9 ? 3'h3 : _GEN_110; // @[Conditional.scala 39:67 PEArray.scala 132:19]
  wire [2:0] _GEN_112 = _T_8 ? 3'h2 : _GEN_111; // @[Conditional.scala 39:67 PEArray.scala 128:19]
  wire [2:0] _GEN_113 = _T_7 ? 3'h1 : _GEN_112; // @[Conditional.scala 39:67 PEArray.scala 124:19]
  wire [7:0] _GEN_118 = io_control_signal_mask[4] ? io_control_signal_gru_out_width : {{2'd0}, GRU_out_width}; // @[PEArray.scala 116:57 PEArray.scala 145:23 PEArray.scala 104:26]
  wire [9:0] _count_T_1 = count + 10'h1; // @[PEArray.scala 162:24]
  wire [9:0] _GEN_120 = count != 10'h33 ? _count_T_1 : count; // @[PEArray.scala 161:27 PEArray.scala 162:15 PEArray.scala 101:22]
  wire [9:0] _GEN_124 = count != 10'h188 ? _count_T_1 : count; // @[PEArray.scala 183:28 PEArray.scala 184:15 PEArray.scala 101:22]
  wire [9:0] _GEN_125 = count == 10'h188 ? 10'h0 : _GEN_124; // @[PEArray.scala 186:28 PEArray.scala 187:15]
  wire [2:0] _GEN_126 = count == 10'h188 ? 3'h0 : state; // @[PEArray.scala 186:28 PEArray.scala 188:15 PEArray.scala 100:22]
  wire [9:0] _GEN_127 = count != count_max ? _count_T_1 : count; // @[PEArray.scala 192:32 PEArray.scala 193:15 PEArray.scala 101:22]
  wire [5:0] _GEN_128 = count == 10'h0 ? L0index_begin : L0Index; // @[PEArray.scala 195:26 PEArray.scala 196:17 PEArray.scala 39:24]
  wire [9:0] _T_27 = count_max - 10'h1; // @[PEArray.scala 198:51]
  wire [15:0] _GEN_129 = 6'h0 == L0Index ? io_FromL1 : L0Memory_0; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_130 = 6'h1 == L0Index ? io_FromL1 : L0Memory_1; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_131 = 6'h2 == L0Index ? io_FromL1 : L0Memory_2; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_132 = 6'h3 == L0Index ? io_FromL1 : L0Memory_3; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_133 = 6'h4 == L0Index ? io_FromL1 : L0Memory_4; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_134 = 6'h5 == L0Index ? io_FromL1 : L0Memory_5; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_135 = 6'h6 == L0Index ? io_FromL1 : L0Memory_6; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_136 = 6'h7 == L0Index ? io_FromL1 : L0Memory_7; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_137 = 6'h8 == L0Index ? io_FromL1 : L0Memory_8; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_138 = 6'h9 == L0Index ? io_FromL1 : L0Memory_9; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_139 = 6'ha == L0Index ? io_FromL1 : L0Memory_10; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_140 = 6'hb == L0Index ? io_FromL1 : L0Memory_11; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_141 = 6'hc == L0Index ? io_FromL1 : L0Memory_12; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_142 = 6'hd == L0Index ? io_FromL1 : L0Memory_13; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_143 = 6'he == L0Index ? io_FromL1 : L0Memory_14; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_144 = 6'hf == L0Index ? io_FromL1 : L0Memory_15; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_145 = 6'h10 == L0Index ? io_FromL1 : L0Memory_16; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_146 = 6'h11 == L0Index ? io_FromL1 : L0Memory_17; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_147 = 6'h12 == L0Index ? io_FromL1 : L0Memory_18; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_148 = 6'h13 == L0Index ? io_FromL1 : L0Memory_19; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_149 = 6'h14 == L0Index ? io_FromL1 : L0Memory_20; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_150 = 6'h15 == L0Index ? io_FromL1 : L0Memory_21; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_151 = 6'h16 == L0Index ? io_FromL1 : L0Memory_22; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_152 = 6'h17 == L0Index ? io_FromL1 : L0Memory_23; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_153 = 6'h18 == L0Index ? io_FromL1 : L0Memory_24; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_154 = 6'h19 == L0Index ? io_FromL1 : L0Memory_25; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_155 = 6'h1a == L0Index ? io_FromL1 : L0Memory_26; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_156 = 6'h1b == L0Index ? io_FromL1 : L0Memory_27; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_157 = 6'h1c == L0Index ? io_FromL1 : L0Memory_28; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_158 = 6'h1d == L0Index ? io_FromL1 : L0Memory_29; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_159 = 6'h1e == L0Index ? io_FromL1 : L0Memory_30; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_160 = 6'h1f == L0Index ? io_FromL1 : L0Memory_31; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_161 = 6'h20 == L0Index ? io_FromL1 : L0Memory_32; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_162 = 6'h21 == L0Index ? io_FromL1 : L0Memory_33; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_163 = 6'h22 == L0Index ? io_FromL1 : L0Memory_34; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_164 = 6'h23 == L0Index ? io_FromL1 : L0Memory_35; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_165 = 6'h24 == L0Index ? io_FromL1 : L0Memory_36; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_166 = 6'h25 == L0Index ? io_FromL1 : L0Memory_37; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_167 = 6'h26 == L0Index ? io_FromL1 : L0Memory_38; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_168 = 6'h27 == L0Index ? io_FromL1 : L0Memory_39; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_169 = 6'h28 == L0Index ? io_FromL1 : L0Memory_40; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_170 = 6'h29 == L0Index ? io_FromL1 : L0Memory_41; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_171 = 6'h2a == L0Index ? io_FromL1 : L0Memory_42; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_172 = 6'h2b == L0Index ? io_FromL1 : L0Memory_43; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_173 = 6'h2c == L0Index ? io_FromL1 : L0Memory_44; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_174 = 6'h2d == L0Index ? io_FromL1 : L0Memory_45; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_175 = 6'h2e == L0Index ? io_FromL1 : L0Memory_46; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_176 = 6'h2f == L0Index ? io_FromL1 : L0Memory_47; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_177 = 6'h30 == L0Index ? io_FromL1 : L0Memory_48; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_178 = 6'h31 == L0Index ? io_FromL1 : L0Memory_49; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_179 = 6'h32 == L0Index ? io_FromL1 : L0Memory_50; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_180 = 6'h33 == L0Index ? io_FromL1 : L0Memory_51; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_181 = 6'h34 == L0Index ? io_FromL1 : L0Memory_52; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_182 = 6'h35 == L0Index ? io_FromL1 : L0Memory_53; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_183 = 6'h36 == L0Index ? io_FromL1 : L0Memory_54; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_184 = 6'h37 == L0Index ? io_FromL1 : L0Memory_55; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_185 = 6'h38 == L0Index ? io_FromL1 : L0Memory_56; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_186 = 6'h39 == L0Index ? io_FromL1 : L0Memory_57; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_187 = 6'h3a == L0Index ? io_FromL1 : L0Memory_58; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_188 = 6'h3b == L0Index ? io_FromL1 : L0Memory_59; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_189 = 6'h3c == L0Index ? io_FromL1 : L0Memory_60; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_190 = 6'h3d == L0Index ? io_FromL1 : L0Memory_61; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_191 = 6'h3e == L0Index ? io_FromL1 : L0Memory_62; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_192 = 6'h3f == L0Index ? io_FromL1 : L0Memory_63; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_193 = 7'h40 == _GEN_793 ? io_FromL1 : L0Memory_64; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_194 = 7'h41 == _GEN_793 ? io_FromL1 : L0Memory_65; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_195 = 7'h42 == _GEN_793 ? io_FromL1 : L0Memory_66; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_196 = 7'h43 == _GEN_793 ? io_FromL1 : L0Memory_67; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_197 = 7'h44 == _GEN_793 ? io_FromL1 : L0Memory_68; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_198 = 7'h45 == _GEN_793 ? io_FromL1 : L0Memory_69; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_199 = 7'h46 == _GEN_793 ? io_FromL1 : L0Memory_70; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_200 = 7'h47 == _GEN_793 ? io_FromL1 : L0Memory_71; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_201 = 7'h48 == _GEN_793 ? io_FromL1 : L0Memory_72; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_202 = 7'h49 == _GEN_793 ? io_FromL1 : L0Memory_73; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_203 = 7'h4a == _GEN_793 ? io_FromL1 : L0Memory_74; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_204 = 7'h4b == _GEN_793 ? io_FromL1 : L0Memory_75; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_205 = 7'h4c == _GEN_793 ? io_FromL1 : L0Memory_76; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_206 = 7'h4d == _GEN_793 ? io_FromL1 : L0Memory_77; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_207 = 7'h4e == _GEN_793 ? io_FromL1 : L0Memory_78; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_208 = 7'h4f == _GEN_793 ? io_FromL1 : L0Memory_79; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_209 = 7'h50 == _GEN_793 ? io_FromL1 : L0Memory_80; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_210 = 7'h51 == _GEN_793 ? io_FromL1 : L0Memory_81; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_211 = 7'h52 == _GEN_793 ? io_FromL1 : L0Memory_82; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_212 = 7'h53 == _GEN_793 ? io_FromL1 : L0Memory_83; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_213 = 7'h54 == _GEN_793 ? io_FromL1 : L0Memory_84; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_214 = 7'h55 == _GEN_793 ? io_FromL1 : L0Memory_85; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_215 = 7'h56 == _GEN_793 ? io_FromL1 : L0Memory_86; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_216 = 7'h57 == _GEN_793 ? io_FromL1 : L0Memory_87; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_217 = 7'h58 == _GEN_793 ? io_FromL1 : L0Memory_88; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_218 = 7'h59 == _GEN_793 ? io_FromL1 : L0Memory_89; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_219 = 7'h5a == _GEN_793 ? io_FromL1 : L0Memory_90; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_220 = 7'h5b == _GEN_793 ? io_FromL1 : L0Memory_91; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_221 = 7'h5c == _GEN_793 ? io_FromL1 : L0Memory_92; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_222 = 7'h5d == _GEN_793 ? io_FromL1 : L0Memory_93; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_223 = 7'h5e == _GEN_793 ? io_FromL1 : L0Memory_94; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_224 = 7'h5f == _GEN_793 ? io_FromL1 : L0Memory_95; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_225 = 7'h60 == _GEN_793 ? io_FromL1 : L0Memory_96; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_226 = 7'h61 == _GEN_793 ? io_FromL1 : L0Memory_97; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_227 = 7'h62 == _GEN_793 ? io_FromL1 : L0Memory_98; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_228 = 7'h63 == _GEN_793 ? io_FromL1 : L0Memory_99; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [5:0] _L0Index_T_2 = L0Index + 6'h1; // @[PEArray.scala 200:28]
  wire [15:0] _GEN_229 = count >= 10'h1 & count <= _T_27 ? _GEN_129 : L0Memory_0; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_230 = count >= 10'h1 & count <= _T_27 ? _GEN_130 : L0Memory_1; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_231 = count >= 10'h1 & count <= _T_27 ? _GEN_131 : L0Memory_2; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_232 = count >= 10'h1 & count <= _T_27 ? _GEN_132 : L0Memory_3; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_233 = count >= 10'h1 & count <= _T_27 ? _GEN_133 : L0Memory_4; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_234 = count >= 10'h1 & count <= _T_27 ? _GEN_134 : L0Memory_5; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_235 = count >= 10'h1 & count <= _T_27 ? _GEN_135 : L0Memory_6; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_236 = count >= 10'h1 & count <= _T_27 ? _GEN_136 : L0Memory_7; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_237 = count >= 10'h1 & count <= _T_27 ? _GEN_137 : L0Memory_8; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_238 = count >= 10'h1 & count <= _T_27 ? _GEN_138 : L0Memory_9; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_239 = count >= 10'h1 & count <= _T_27 ? _GEN_139 : L0Memory_10; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_240 = count >= 10'h1 & count <= _T_27 ? _GEN_140 : L0Memory_11; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_241 = count >= 10'h1 & count <= _T_27 ? _GEN_141 : L0Memory_12; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_242 = count >= 10'h1 & count <= _T_27 ? _GEN_142 : L0Memory_13; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_243 = count >= 10'h1 & count <= _T_27 ? _GEN_143 : L0Memory_14; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_244 = count >= 10'h1 & count <= _T_27 ? _GEN_144 : L0Memory_15; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_245 = count >= 10'h1 & count <= _T_27 ? _GEN_145 : L0Memory_16; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_246 = count >= 10'h1 & count <= _T_27 ? _GEN_146 : L0Memory_17; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_247 = count >= 10'h1 & count <= _T_27 ? _GEN_147 : L0Memory_18; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_248 = count >= 10'h1 & count <= _T_27 ? _GEN_148 : L0Memory_19; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_249 = count >= 10'h1 & count <= _T_27 ? _GEN_149 : L0Memory_20; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_250 = count >= 10'h1 & count <= _T_27 ? _GEN_150 : L0Memory_21; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_251 = count >= 10'h1 & count <= _T_27 ? _GEN_151 : L0Memory_22; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_252 = count >= 10'h1 & count <= _T_27 ? _GEN_152 : L0Memory_23; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_253 = count >= 10'h1 & count <= _T_27 ? _GEN_153 : L0Memory_24; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_254 = count >= 10'h1 & count <= _T_27 ? _GEN_154 : L0Memory_25; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_255 = count >= 10'h1 & count <= _T_27 ? _GEN_155 : L0Memory_26; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_256 = count >= 10'h1 & count <= _T_27 ? _GEN_156 : L0Memory_27; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_257 = count >= 10'h1 & count <= _T_27 ? _GEN_157 : L0Memory_28; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_258 = count >= 10'h1 & count <= _T_27 ? _GEN_158 : L0Memory_29; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_259 = count >= 10'h1 & count <= _T_27 ? _GEN_159 : L0Memory_30; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_260 = count >= 10'h1 & count <= _T_27 ? _GEN_160 : L0Memory_31; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_261 = count >= 10'h1 & count <= _T_27 ? _GEN_161 : L0Memory_32; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_262 = count >= 10'h1 & count <= _T_27 ? _GEN_162 : L0Memory_33; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_263 = count >= 10'h1 & count <= _T_27 ? _GEN_163 : L0Memory_34; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_264 = count >= 10'h1 & count <= _T_27 ? _GEN_164 : L0Memory_35; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_265 = count >= 10'h1 & count <= _T_27 ? _GEN_165 : L0Memory_36; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_266 = count >= 10'h1 & count <= _T_27 ? _GEN_166 : L0Memory_37; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_267 = count >= 10'h1 & count <= _T_27 ? _GEN_167 : L0Memory_38; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_268 = count >= 10'h1 & count <= _T_27 ? _GEN_168 : L0Memory_39; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_269 = count >= 10'h1 & count <= _T_27 ? _GEN_169 : L0Memory_40; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_270 = count >= 10'h1 & count <= _T_27 ? _GEN_170 : L0Memory_41; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_271 = count >= 10'h1 & count <= _T_27 ? _GEN_171 : L0Memory_42; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_272 = count >= 10'h1 & count <= _T_27 ? _GEN_172 : L0Memory_43; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_273 = count >= 10'h1 & count <= _T_27 ? _GEN_173 : L0Memory_44; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_274 = count >= 10'h1 & count <= _T_27 ? _GEN_174 : L0Memory_45; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_275 = count >= 10'h1 & count <= _T_27 ? _GEN_175 : L0Memory_46; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_276 = count >= 10'h1 & count <= _T_27 ? _GEN_176 : L0Memory_47; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_277 = count >= 10'h1 & count <= _T_27 ? _GEN_177 : L0Memory_48; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_278 = count >= 10'h1 & count <= _T_27 ? _GEN_178 : L0Memory_49; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_279 = count >= 10'h1 & count <= _T_27 ? _GEN_179 : L0Memory_50; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_280 = count >= 10'h1 & count <= _T_27 ? _GEN_180 : L0Memory_51; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_281 = count >= 10'h1 & count <= _T_27 ? _GEN_181 : L0Memory_52; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_282 = count >= 10'h1 & count <= _T_27 ? _GEN_182 : L0Memory_53; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_283 = count >= 10'h1 & count <= _T_27 ? _GEN_183 : L0Memory_54; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_284 = count >= 10'h1 & count <= _T_27 ? _GEN_184 : L0Memory_55; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_285 = count >= 10'h1 & count <= _T_27 ? _GEN_185 : L0Memory_56; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_286 = count >= 10'h1 & count <= _T_27 ? _GEN_186 : L0Memory_57; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_287 = count >= 10'h1 & count <= _T_27 ? _GEN_187 : L0Memory_58; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_288 = count >= 10'h1 & count <= _T_27 ? _GEN_188 : L0Memory_59; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_289 = count >= 10'h1 & count <= _T_27 ? _GEN_189 : L0Memory_60; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_290 = count >= 10'h1 & count <= _T_27 ? _GEN_190 : L0Memory_61; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_291 = count >= 10'h1 & count <= _T_27 ? _GEN_191 : L0Memory_62; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_292 = count >= 10'h1 & count <= _T_27 ? _GEN_192 : L0Memory_63; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_293 = count >= 10'h1 & count <= _T_27 ? _GEN_193 : L0Memory_64; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_294 = count >= 10'h1 & count <= _T_27 ? _GEN_194 : L0Memory_65; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_295 = count >= 10'h1 & count <= _T_27 ? _GEN_195 : L0Memory_66; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_296 = count >= 10'h1 & count <= _T_27 ? _GEN_196 : L0Memory_67; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_297 = count >= 10'h1 & count <= _T_27 ? _GEN_197 : L0Memory_68; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_298 = count >= 10'h1 & count <= _T_27 ? _GEN_198 : L0Memory_69; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_299 = count >= 10'h1 & count <= _T_27 ? _GEN_199 : L0Memory_70; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_300 = count >= 10'h1 & count <= _T_27 ? _GEN_200 : L0Memory_71; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_301 = count >= 10'h1 & count <= _T_27 ? _GEN_201 : L0Memory_72; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_302 = count >= 10'h1 & count <= _T_27 ? _GEN_202 : L0Memory_73; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_303 = count >= 10'h1 & count <= _T_27 ? _GEN_203 : L0Memory_74; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_304 = count >= 10'h1 & count <= _T_27 ? _GEN_204 : L0Memory_75; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_305 = count >= 10'h1 & count <= _T_27 ? _GEN_205 : L0Memory_76; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_306 = count >= 10'h1 & count <= _T_27 ? _GEN_206 : L0Memory_77; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_307 = count >= 10'h1 & count <= _T_27 ? _GEN_207 : L0Memory_78; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_308 = count >= 10'h1 & count <= _T_27 ? _GEN_208 : L0Memory_79; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_309 = count >= 10'h1 & count <= _T_27 ? _GEN_209 : L0Memory_80; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_310 = count >= 10'h1 & count <= _T_27 ? _GEN_210 : L0Memory_81; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_311 = count >= 10'h1 & count <= _T_27 ? _GEN_211 : L0Memory_82; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_312 = count >= 10'h1 & count <= _T_27 ? _GEN_212 : L0Memory_83; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_313 = count >= 10'h1 & count <= _T_27 ? _GEN_213 : L0Memory_84; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_314 = count >= 10'h1 & count <= _T_27 ? _GEN_214 : L0Memory_85; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_315 = count >= 10'h1 & count <= _T_27 ? _GEN_215 : L0Memory_86; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_316 = count >= 10'h1 & count <= _T_27 ? _GEN_216 : L0Memory_87; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_317 = count >= 10'h1 & count <= _T_27 ? _GEN_217 : L0Memory_88; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_318 = count >= 10'h1 & count <= _T_27 ? _GEN_218 : L0Memory_89; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_319 = count >= 10'h1 & count <= _T_27 ? _GEN_219 : L0Memory_90; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_320 = count >= 10'h1 & count <= _T_27 ? _GEN_220 : L0Memory_91; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_321 = count >= 10'h1 & count <= _T_27 ? _GEN_221 : L0Memory_92; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_322 = count >= 10'h1 & count <= _T_27 ? _GEN_222 : L0Memory_93; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_323 = count >= 10'h1 & count <= _T_27 ? _GEN_223 : L0Memory_94; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_324 = count >= 10'h1 & count <= _T_27 ? _GEN_224 : L0Memory_95; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_325 = count >= 10'h1 & count <= _T_27 ? _GEN_225 : L0Memory_96; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_326 = count >= 10'h1 & count <= _T_27 ? _GEN_226 : L0Memory_97; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_327 = count >= 10'h1 & count <= _T_27 ? _GEN_227 : L0Memory_98; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_328 = count >= 10'h1 & count <= _T_27 ? _GEN_228 : L0Memory_99; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [5:0] _GEN_329 = count >= 10'h1 & count <= _T_27 ? _L0Index_T_2 : _GEN_128; // @[PEArray.scala 198:59 PEArray.scala 200:17]
  wire [9:0] _GEN_330 = count == count_max ? 10'h0 : _GEN_127; // @[PEArray.scala 202:32 PEArray.scala 203:15]
  wire [2:0] _GEN_331 = count == count_max ? 3'h0 : state; // @[PEArray.scala 202:32 PEArray.scala 204:15 PEArray.scala 100:22]
  wire [9:0] _GEN_865 = {{4'd0}, GRU_out_width}; // @[PEArray.scala 220:19]
  wire [9:0] _GEN_0 = count % _GEN_865; // @[PEArray.scala 220:19]
  wire [5:0] _T_36 = _GEN_0[5:0]; // @[PEArray.scala 220:19]
  wire [5:0] _T_38 = GRU_out_width - 6'h1; // @[PEArray.scala 220:55]
  wire [5:0] _GEN_334 = _T_36 == _T_38 ? _L0Index_T_2 : L0index_begin; // @[PEArray.scala 220:62 PEArray.scala 221:17 PEArray.scala 214:15]
  wire [5:0] _GEN_346 = _T_41 ? _GEN_334 : L0Index; // @[Conditional.scala 39:67 PEArray.scala 39:24]
  wire [9:0] _GEN_347 = _T_41 ? _GEN_330 : count; // @[Conditional.scala 39:67 PEArray.scala 101:22]
  wire [2:0] _GEN_348 = _T_41 ? _GEN_331 : state; // @[Conditional.scala 39:67 PEArray.scala 100:22]
  wire [5:0] _GEN_353 = _T_31 ? _GEN_334 : _GEN_346; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_354 = _T_31 ? _GEN_330 : _GEN_347; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_355 = _T_31 ? _GEN_331 : _GEN_348; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_356 = _T_22 ? _GEN_330 : _GEN_354; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_357 = _T_22 ? _GEN_329 : _GEN_353; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_458 = _T_22 ? _GEN_331 : _GEN_355; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_690 = _T_3 ? _GEN_118 : {{2'd0}, GRU_out_width}; // @[Conditional.scala 40:58 PEArray.scala 104:26]
  FP16MulAdder FP16MAC ( // @[PEArray.scala 72:23]
    .io_a(FP16MAC_io_a),
    .io_b(FP16MAC_io_b),
    .io_c(FP16MAC_io_c),
    .io_out(FP16MAC_io_out)
  );
  assign io_ToRightPE = mux3out_reg; // @[PEArray.scala 95:16]
  assign io_ToBelowPE = mux2out_reg; // @[PEArray.scala 94:16]
  assign FP16MAC_io_a = sel1 ? io_FromL1 : io_FromLeftPE; // @[PEArray.scala 50:14 PEArray.scala 50:23 PEArray.scala 51:24]
  assign FP16MAC_io_b = sel5 ? mux4out : _GEN_105; // @[PEArray.scala 77:13 PEArray.scala 78:18 PEArray.scala 81:18]
  assign FP16MAC_io_c = sel5 ? _GEN_105 : mux4out; // @[PEArray.scala 77:13 PEArray.scala 79:18 PEArray.scala 82:18]
  always @(posedge clock) begin
    if (reset) begin // @[PEArray.scala 39:24]
      L0Index <= 6'h0; // @[PEArray.scala 39:24]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h2; // @[PEArray.scala 159:15]
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        L0Index <= 6'ha; // @[PEArray.scala 181:15]
      end else begin
        L0Index <= _GEN_357;
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_0 <= _GEN_229;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_1 <= _GEN_230;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_2 <= _GEN_231;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_3 <= _GEN_232;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_4 <= _GEN_233;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_5 <= _GEN_234;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_6 <= _GEN_235;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_7 <= _GEN_236;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_8 <= _GEN_237;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_9 <= _GEN_238;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_10 <= _GEN_239;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_11 <= _GEN_240;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_12 <= _GEN_241;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_13 <= _GEN_242;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_14 <= _GEN_243;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_15 <= _GEN_244;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_16 <= _GEN_245;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_17 <= _GEN_246;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_18 <= _GEN_247;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_19 <= _GEN_248;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_20 <= _GEN_249;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_21 <= _GEN_250;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_22 <= _GEN_251;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_23 <= _GEN_252;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_24 <= _GEN_253;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_25 <= _GEN_254;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_26 <= _GEN_255;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_27 <= _GEN_256;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_28 <= _GEN_257;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_29 <= _GEN_258;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_30 <= _GEN_259;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_31 <= _GEN_260;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_32 <= _GEN_261;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_33 <= _GEN_262;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_34 <= _GEN_263;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_35 <= _GEN_264;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_36 <= _GEN_265;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_37 <= _GEN_266;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_38 <= _GEN_267;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_39 <= _GEN_268;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_40 <= _GEN_269;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_41 <= _GEN_270;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_42 <= _GEN_271;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_43 <= _GEN_272;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_44 <= _GEN_273;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_45 <= _GEN_274;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_46 <= _GEN_275;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_47 <= _GEN_276;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_48 <= _GEN_277;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_49 <= _GEN_278;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_50 <= _GEN_279;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_51 <= _GEN_280;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_52 <= _GEN_281;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_53 <= _GEN_282;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_54 <= _GEN_283;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_55 <= _GEN_284;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_56 <= _GEN_285;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_57 <= _GEN_286;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_58 <= _GEN_287;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_59 <= _GEN_288;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_60 <= _GEN_289;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_61 <= _GEN_290;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_62 <= _GEN_291;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_63 <= _GEN_292;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_64 <= _GEN_293;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_65 <= _GEN_294;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_66 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_67 <= _GEN_296;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_68 <= _GEN_297;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_69 <= _GEN_298;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_70 <= _GEN_299;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_71 <= _GEN_300;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_72 <= _GEN_301;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_73 <= _GEN_302;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_74 <= _GEN_303;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_75 <= _GEN_304;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_76 <= _GEN_305;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_77 <= _GEN_306;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_78 <= _GEN_307;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_79 <= _GEN_308;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_80 <= _GEN_309;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_81 <= _GEN_310;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_82 <= _GEN_311;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_83 <= _GEN_312;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_84 <= _GEN_313;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_85 <= _GEN_314;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_86 <= _GEN_315;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_87 <= _GEN_316;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_88 <= _GEN_317;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_89 <= _GEN_318;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_90 <= _GEN_319;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_91 <= _GEN_320;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_92 <= _GEN_321;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_93 <= _GEN_322;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_94 <= _GEN_323;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_95 <= _GEN_324;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_96 <= _GEN_325;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_97 <= _GEN_326;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_98 <= _GEN_327;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_99 <= _GEN_328;
          end
        end
      end
    end
    if (reset) begin // @[PEArray.scala 100:22]
      state <= 3'h0; // @[PEArray.scala 100:22]
    end else if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[4]) begin // @[PEArray.scala 116:57]
        if (_T_6) begin // @[Conditional.scala 40:58]
          state <= 3'h0; // @[PEArray.scala 120:19]
        end else begin
          state <= _GEN_113;
        end
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      if (count == 10'h33) begin // @[PEArray.scala 164:27]
        state <= 3'h0; // @[PEArray.scala 166:15]
      end
    end else if (_T_16) begin // @[Conditional.scala 39:67]
      state <= _GEN_126;
    end else begin
      state <= _GEN_458;
    end
    if (reset) begin // @[PEArray.scala 90:28]
      mux2out_reg <= 16'h0; // @[PEArray.scala 90:28]
    end else begin
      mux2out_reg <= MAC_out; // @[PEArray.scala 90:28]
    end
    if (reset) begin // @[PEArray.scala 91:28]
      mux3out_reg <= 16'h0; // @[PEArray.scala 91:28]
    end else if (sel3) begin // @[PEArray.scala 56:14]
      mux3out_reg <= MAC_out; // @[PEArray.scala 56:23]
    end else if (sel1) begin // @[PEArray.scala 50:14]
      mux3out_reg <= io_FromL1; // @[PEArray.scala 50:23]
    end else begin
      mux3out_reg <= io_FromLeftPE; // @[PEArray.scala 51:24]
    end
    if (reset) begin // @[PEArray.scala 101:22]
      count <= 10'h0; // @[PEArray.scala 101:22]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        if (count == 10'h33) begin // @[PEArray.scala 164:27]
          count <= 10'h0; // @[PEArray.scala 165:15]
        end else begin
          count <= _GEN_120;
        end
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        count <= _GEN_125;
      end else begin
        count <= _GEN_356;
      end
    end
    if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[4]) begin // @[PEArray.scala 116:57]
        count_max <= io_control_signal_count; // @[PEArray.scala 143:19]
      end
    end
    if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[4]) begin // @[PEArray.scala 116:57]
        L0index_begin <= io_control_signal_L0index; // @[PEArray.scala 144:23]
      end
    end
    GRU_out_width <= _GEN_690[5:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  L0Index = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  L0Memory_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  L0Memory_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  L0Memory_2 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  L0Memory_3 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  L0Memory_4 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  L0Memory_5 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  L0Memory_6 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  L0Memory_7 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  L0Memory_8 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  L0Memory_9 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  L0Memory_10 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  L0Memory_11 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  L0Memory_12 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  L0Memory_13 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  L0Memory_14 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  L0Memory_15 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  L0Memory_16 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  L0Memory_17 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  L0Memory_18 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  L0Memory_19 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  L0Memory_20 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  L0Memory_21 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  L0Memory_22 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  L0Memory_23 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  L0Memory_24 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  L0Memory_25 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  L0Memory_26 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  L0Memory_27 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  L0Memory_28 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  L0Memory_29 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  L0Memory_30 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  L0Memory_31 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  L0Memory_32 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  L0Memory_33 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  L0Memory_34 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  L0Memory_35 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  L0Memory_36 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  L0Memory_37 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  L0Memory_38 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  L0Memory_39 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  L0Memory_40 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  L0Memory_41 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  L0Memory_42 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  L0Memory_43 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  L0Memory_44 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  L0Memory_45 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  L0Memory_46 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  L0Memory_47 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  L0Memory_48 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  L0Memory_49 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  L0Memory_50 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  L0Memory_51 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  L0Memory_52 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  L0Memory_53 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  L0Memory_54 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  L0Memory_55 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  L0Memory_56 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  L0Memory_57 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  L0Memory_58 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  L0Memory_59 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  L0Memory_60 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  L0Memory_61 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  L0Memory_62 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  L0Memory_63 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  L0Memory_64 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  L0Memory_65 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  L0Memory_66 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  L0Memory_67 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  L0Memory_68 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  L0Memory_69 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  L0Memory_70 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  L0Memory_71 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  L0Memory_72 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  L0Memory_73 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  L0Memory_74 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  L0Memory_75 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  L0Memory_76 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  L0Memory_77 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  L0Memory_78 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  L0Memory_79 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  L0Memory_80 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  L0Memory_81 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  L0Memory_82 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  L0Memory_83 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  L0Memory_84 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  L0Memory_85 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  L0Memory_86 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  L0Memory_87 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  L0Memory_88 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  L0Memory_89 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  L0Memory_90 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  L0Memory_91 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  L0Memory_92 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  L0Memory_93 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  L0Memory_94 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  L0Memory_95 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  L0Memory_96 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  L0Memory_97 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  L0Memory_98 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  L0Memory_99 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  state = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  mux2out_reg = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  mux3out_reg = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  count = _RAND_104[9:0];
  _RAND_105 = {1{`RANDOM}};
  count_max = _RAND_105[9:0];
  _RAND_106 = {1{`RANDOM}};
  L0index_begin = _RAND_106[5:0];
  _RAND_107 = {1{`RANDOM}};
  GRU_out_width = _RAND_107[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PE_24(
  input         clock,
  input         reset,
  input  [15:0] io_FromAbovePE,
  input  [15:0] io_FromLeftPE,
  input  [15:0] io_FromL1,
  input  [11:0] io_control_signal_mask,
  output [15:0] io_ToRightPE,
  output [15:0] io_ToBelowPE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] FP16MAC_io_a; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_b; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_c; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_out; // @[PEArray.scala 72:23]
  reg [5:0] L0Index; // @[PEArray.scala 39:24]
  reg [15:0] L0Memory_0; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_1; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_2; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_3; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_4; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_5; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_6; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_7; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_8; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_9; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_10; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_11; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_12; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_13; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_14; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_15; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_16; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_17; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_18; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_19; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_20; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_21; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_22; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_23; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_24; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_25; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_26; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_27; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_28; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_29; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_30; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_31; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_32; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_33; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_34; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_35; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_36; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_37; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_38; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_39; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_40; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_41; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_42; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_43; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_44; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_45; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_46; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_47; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_48; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_49; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_50; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_51; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_52; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_53; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_54; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_55; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_56; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_57; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_58; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_59; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_60; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_61; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_62; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_63; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_64; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_65; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_66; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_67; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_68; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_69; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_70; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_71; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_72; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_73; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_74; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_75; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_76; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_77; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_78; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_79; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_80; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_81; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_82; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_83; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_84; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_85; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_86; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_87; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_88; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_89; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_90; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_91; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_92; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_93; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_94; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_95; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_96; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_97; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_98; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_99; // @[PEArray.scala 40:21]
  reg [2:0] state; // @[PEArray.scala 100:22]
  wire  _T_3 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_12 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_16 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_22 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_31 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_41 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_342 = _T_41 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 231:12 PEArray.scala 32:8]
  wire  _GEN_349 = _T_31 ? 1'h0 : _GEN_342; // @[Conditional.scala 39:67 PEArray.scala 208:12]
  wire  _GEN_459 = _T_22 | _GEN_349; // @[Conditional.scala 39:67 PEArray.scala 32:8]
  wire  _GEN_463 = _T_16 ? 1'h0 : _GEN_459; // @[Conditional.scala 39:67]
  wire  _GEN_572 = _T_12 | _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 149:12]
  wire  sel1 = _T_3 | _GEN_572; // @[Conditional.scala 40:58 PEArray.scala 108:12]
  wire [15:0] MAC_out = FP16MAC_io_out; // @[PEArray.scala 47:21 PEArray.scala 85:11]
  wire  _GEN_465 = _T_16 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 177:12]
  wire  _GEN_580 = _T_12 | _GEN_465; // @[Conditional.scala 39:67 PEArray.scala 34:8]
  wire  sel3 = _T_3 | _GEN_580; // @[Conditional.scala 40:58 PEArray.scala 110:12]
  wire [1:0] _GEN_344 = _T_41 ? 2'h2 : 2'h0; // @[Conditional.scala 39:67 PEArray.scala 233:12 PEArray.scala 35:8]
  wire [1:0] _GEN_351 = _T_31 ? 2'h2 : _GEN_344; // @[Conditional.scala 39:67 PEArray.scala 210:12]
  wire [1:0] _GEN_461 = _T_22 ? 2'h0 : _GEN_351; // @[Conditional.scala 39:67 PEArray.scala 35:8]
  wire [1:0] _GEN_466 = _T_16 ? 2'h0 : _GEN_461; // @[Conditional.scala 39:67 PEArray.scala 178:12]
  wire [1:0] _GEN_574 = _T_12 ? 2'h0 : _GEN_466; // @[Conditional.scala 39:67]
  wire [1:0] sel4 = _T_3 ? 2'h0 : _GEN_574; // @[Conditional.scala 40:58 PEArray.scala 111:12]
  wire [15:0] _GEN_3 = sel4 == 2'h2 ? io_FromL1 : 16'h0; // @[PEArray.scala 65:28 PEArray.scala 66:15 PEArray.scala 69:15]
  wire [15:0] _GEN_4 = sel4 == 2'h1 ? io_FromAbovePE : _GEN_3; // @[PEArray.scala 62:28 PEArray.scala 63:15]
  wire [15:0] mux4out = sel4 == 2'h0 ? 16'h0 : _GEN_4; // @[PEArray.scala 59:22 PEArray.scala 60:13]
  wire [15:0] _GEN_7 = 6'h1 == L0Index ? L0Memory_1 : L0Memory_0; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_8 = 6'h2 == L0Index ? L0Memory_2 : _GEN_7; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_9 = 6'h3 == L0Index ? L0Memory_3 : _GEN_8; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_10 = 6'h4 == L0Index ? L0Memory_4 : _GEN_9; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_11 = 6'h5 == L0Index ? L0Memory_5 : _GEN_10; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_12 = 6'h6 == L0Index ? L0Memory_6 : _GEN_11; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_13 = 6'h7 == L0Index ? L0Memory_7 : _GEN_12; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_14 = 6'h8 == L0Index ? L0Memory_8 : _GEN_13; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_15 = 6'h9 == L0Index ? L0Memory_9 : _GEN_14; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_16 = 6'ha == L0Index ? L0Memory_10 : _GEN_15; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_17 = 6'hb == L0Index ? L0Memory_11 : _GEN_16; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_18 = 6'hc == L0Index ? L0Memory_12 : _GEN_17; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_19 = 6'hd == L0Index ? L0Memory_13 : _GEN_18; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_20 = 6'he == L0Index ? L0Memory_14 : _GEN_19; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_21 = 6'hf == L0Index ? L0Memory_15 : _GEN_20; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_22 = 6'h10 == L0Index ? L0Memory_16 : _GEN_21; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_23 = 6'h11 == L0Index ? L0Memory_17 : _GEN_22; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_24 = 6'h12 == L0Index ? L0Memory_18 : _GEN_23; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_25 = 6'h13 == L0Index ? L0Memory_19 : _GEN_24; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_26 = 6'h14 == L0Index ? L0Memory_20 : _GEN_25; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_27 = 6'h15 == L0Index ? L0Memory_21 : _GEN_26; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_28 = 6'h16 == L0Index ? L0Memory_22 : _GEN_27; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_29 = 6'h17 == L0Index ? L0Memory_23 : _GEN_28; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_30 = 6'h18 == L0Index ? L0Memory_24 : _GEN_29; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_31 = 6'h19 == L0Index ? L0Memory_25 : _GEN_30; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_32 = 6'h1a == L0Index ? L0Memory_26 : _GEN_31; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_33 = 6'h1b == L0Index ? L0Memory_27 : _GEN_32; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_34 = 6'h1c == L0Index ? L0Memory_28 : _GEN_33; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_35 = 6'h1d == L0Index ? L0Memory_29 : _GEN_34; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_36 = 6'h1e == L0Index ? L0Memory_30 : _GEN_35; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_37 = 6'h1f == L0Index ? L0Memory_31 : _GEN_36; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_38 = 6'h20 == L0Index ? L0Memory_32 : _GEN_37; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_39 = 6'h21 == L0Index ? L0Memory_33 : _GEN_38; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_40 = 6'h22 == L0Index ? L0Memory_34 : _GEN_39; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_41 = 6'h23 == L0Index ? L0Memory_35 : _GEN_40; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_42 = 6'h24 == L0Index ? L0Memory_36 : _GEN_41; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_43 = 6'h25 == L0Index ? L0Memory_37 : _GEN_42; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_44 = 6'h26 == L0Index ? L0Memory_38 : _GEN_43; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_45 = 6'h27 == L0Index ? L0Memory_39 : _GEN_44; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_46 = 6'h28 == L0Index ? L0Memory_40 : _GEN_45; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_47 = 6'h29 == L0Index ? L0Memory_41 : _GEN_46; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_48 = 6'h2a == L0Index ? L0Memory_42 : _GEN_47; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_49 = 6'h2b == L0Index ? L0Memory_43 : _GEN_48; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_50 = 6'h2c == L0Index ? L0Memory_44 : _GEN_49; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_51 = 6'h2d == L0Index ? L0Memory_45 : _GEN_50; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_52 = 6'h2e == L0Index ? L0Memory_46 : _GEN_51; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_53 = 6'h2f == L0Index ? L0Memory_47 : _GEN_52; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_54 = 6'h30 == L0Index ? L0Memory_48 : _GEN_53; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_55 = 6'h31 == L0Index ? L0Memory_49 : _GEN_54; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_56 = 6'h32 == L0Index ? L0Memory_50 : _GEN_55; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_57 = 6'h33 == L0Index ? L0Memory_51 : _GEN_56; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_58 = 6'h34 == L0Index ? L0Memory_52 : _GEN_57; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_59 = 6'h35 == L0Index ? L0Memory_53 : _GEN_58; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_60 = 6'h36 == L0Index ? L0Memory_54 : _GEN_59; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_61 = 6'h37 == L0Index ? L0Memory_55 : _GEN_60; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_62 = 6'h38 == L0Index ? L0Memory_56 : _GEN_61; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_63 = 6'h39 == L0Index ? L0Memory_57 : _GEN_62; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_64 = 6'h3a == L0Index ? L0Memory_58 : _GEN_63; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_65 = 6'h3b == L0Index ? L0Memory_59 : _GEN_64; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_66 = 6'h3c == L0Index ? L0Memory_60 : _GEN_65; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_67 = 6'h3d == L0Index ? L0Memory_61 : _GEN_66; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_68 = 6'h3e == L0Index ? L0Memory_62 : _GEN_67; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_69 = 6'h3f == L0Index ? L0Memory_63 : _GEN_68; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [6:0] _GEN_793 = {{1'd0}, L0Index}; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_70 = 7'h40 == _GEN_793 ? L0Memory_64 : _GEN_69; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_71 = 7'h41 == _GEN_793 ? L0Memory_65 : _GEN_70; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_72 = 7'h42 == _GEN_793 ? L0Memory_66 : _GEN_71; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_73 = 7'h43 == _GEN_793 ? L0Memory_67 : _GEN_72; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_74 = 7'h44 == _GEN_793 ? L0Memory_68 : _GEN_73; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_75 = 7'h45 == _GEN_793 ? L0Memory_69 : _GEN_74; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_76 = 7'h46 == _GEN_793 ? L0Memory_70 : _GEN_75; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_77 = 7'h47 == _GEN_793 ? L0Memory_71 : _GEN_76; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_78 = 7'h48 == _GEN_793 ? L0Memory_72 : _GEN_77; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_79 = 7'h49 == _GEN_793 ? L0Memory_73 : _GEN_78; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_80 = 7'h4a == _GEN_793 ? L0Memory_74 : _GEN_79; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_81 = 7'h4b == _GEN_793 ? L0Memory_75 : _GEN_80; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_82 = 7'h4c == _GEN_793 ? L0Memory_76 : _GEN_81; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_83 = 7'h4d == _GEN_793 ? L0Memory_77 : _GEN_82; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_84 = 7'h4e == _GEN_793 ? L0Memory_78 : _GEN_83; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_85 = 7'h4f == _GEN_793 ? L0Memory_79 : _GEN_84; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_86 = 7'h50 == _GEN_793 ? L0Memory_80 : _GEN_85; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_87 = 7'h51 == _GEN_793 ? L0Memory_81 : _GEN_86; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_88 = 7'h52 == _GEN_793 ? L0Memory_82 : _GEN_87; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_89 = 7'h53 == _GEN_793 ? L0Memory_83 : _GEN_88; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_90 = 7'h54 == _GEN_793 ? L0Memory_84 : _GEN_89; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_91 = 7'h55 == _GEN_793 ? L0Memory_85 : _GEN_90; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_92 = 7'h56 == _GEN_793 ? L0Memory_86 : _GEN_91; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_93 = 7'h57 == _GEN_793 ? L0Memory_87 : _GEN_92; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_94 = 7'h58 == _GEN_793 ? L0Memory_88 : _GEN_93; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_95 = 7'h59 == _GEN_793 ? L0Memory_89 : _GEN_94; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_96 = 7'h5a == _GEN_793 ? L0Memory_90 : _GEN_95; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_97 = 7'h5b == _GEN_793 ? L0Memory_91 : _GEN_96; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_98 = 7'h5c == _GEN_793 ? L0Memory_92 : _GEN_97; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_99 = 7'h5d == _GEN_793 ? L0Memory_93 : _GEN_98; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_100 = 7'h5e == _GEN_793 ? L0Memory_94 : _GEN_99; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_101 = 7'h5f == _GEN_793 ? L0Memory_95 : _GEN_100; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_102 = 7'h60 == _GEN_793 ? L0Memory_96 : _GEN_101; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_103 = 7'h61 == _GEN_793 ? L0Memory_97 : _GEN_102; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_104 = 7'h62 == _GEN_793 ? L0Memory_98 : _GEN_103; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_105 = 7'h63 == _GEN_793 ? L0Memory_99 : _GEN_104; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire  _GEN_575 = _T_12 ? 1'h0 : _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 157:12]
  wire  sel5 = _T_3 ? 1'h0 : _GEN_575; // @[Conditional.scala 40:58 PEArray.scala 112:12]
  reg [15:0] mux2out_reg; // @[PEArray.scala 90:28]
  reg [15:0] mux3out_reg; // @[PEArray.scala 91:28]
  reg [9:0] count; // @[PEArray.scala 101:22]
  reg [5:0] GRU_out_width; // @[PEArray.scala 104:26]
  wire [7:0] _GEN_118 = io_control_signal_mask[3] ? 8'h0 : {{2'd0}, GRU_out_width}; // @[PEArray.scala 116:57 PEArray.scala 145:23 PEArray.scala 104:26]
  wire [9:0] _count_T_1 = count + 10'h1; // @[PEArray.scala 162:24]
  wire [9:0] _GEN_120 = count != 10'h33 ? _count_T_1 : count; // @[PEArray.scala 161:27 PEArray.scala 162:15 PEArray.scala 101:22]
  wire [9:0] _GEN_124 = count != 10'h188 ? _count_T_1 : count; // @[PEArray.scala 183:28 PEArray.scala 184:15 PEArray.scala 101:22]
  wire [9:0] _GEN_125 = count == 10'h188 ? 10'h0 : _GEN_124; // @[PEArray.scala 186:28 PEArray.scala 187:15]
  wire [2:0] _GEN_126 = count == 10'h188 ? 3'h0 : state; // @[PEArray.scala 186:28 PEArray.scala 188:15 PEArray.scala 100:22]
  wire [9:0] _GEN_127 = count != 10'h0 ? _count_T_1 : count; // @[PEArray.scala 192:32 PEArray.scala 193:15 PEArray.scala 101:22]
  wire  _T_24 = count == 10'h0; // @[PEArray.scala 195:18]
  wire [5:0] _GEN_128 = count == 10'h0 ? 6'h0 : L0Index; // @[PEArray.scala 195:26 PEArray.scala 196:17 PEArray.scala 39:24]
  wire [9:0] _T_27 = 10'h0 - 10'h1; // @[PEArray.scala 198:51]
  wire [15:0] _GEN_129 = 6'h0 == L0Index ? io_FromL1 : L0Memory_0; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_130 = 6'h1 == L0Index ? io_FromL1 : L0Memory_1; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_131 = 6'h2 == L0Index ? io_FromL1 : L0Memory_2; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_132 = 6'h3 == L0Index ? io_FromL1 : L0Memory_3; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_133 = 6'h4 == L0Index ? io_FromL1 : L0Memory_4; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_134 = 6'h5 == L0Index ? io_FromL1 : L0Memory_5; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_135 = 6'h6 == L0Index ? io_FromL1 : L0Memory_6; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_136 = 6'h7 == L0Index ? io_FromL1 : L0Memory_7; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_137 = 6'h8 == L0Index ? io_FromL1 : L0Memory_8; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_138 = 6'h9 == L0Index ? io_FromL1 : L0Memory_9; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_139 = 6'ha == L0Index ? io_FromL1 : L0Memory_10; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_140 = 6'hb == L0Index ? io_FromL1 : L0Memory_11; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_141 = 6'hc == L0Index ? io_FromL1 : L0Memory_12; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_142 = 6'hd == L0Index ? io_FromL1 : L0Memory_13; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_143 = 6'he == L0Index ? io_FromL1 : L0Memory_14; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_144 = 6'hf == L0Index ? io_FromL1 : L0Memory_15; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_145 = 6'h10 == L0Index ? io_FromL1 : L0Memory_16; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_146 = 6'h11 == L0Index ? io_FromL1 : L0Memory_17; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_147 = 6'h12 == L0Index ? io_FromL1 : L0Memory_18; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_148 = 6'h13 == L0Index ? io_FromL1 : L0Memory_19; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_149 = 6'h14 == L0Index ? io_FromL1 : L0Memory_20; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_150 = 6'h15 == L0Index ? io_FromL1 : L0Memory_21; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_151 = 6'h16 == L0Index ? io_FromL1 : L0Memory_22; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_152 = 6'h17 == L0Index ? io_FromL1 : L0Memory_23; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_153 = 6'h18 == L0Index ? io_FromL1 : L0Memory_24; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_154 = 6'h19 == L0Index ? io_FromL1 : L0Memory_25; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_155 = 6'h1a == L0Index ? io_FromL1 : L0Memory_26; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_156 = 6'h1b == L0Index ? io_FromL1 : L0Memory_27; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_157 = 6'h1c == L0Index ? io_FromL1 : L0Memory_28; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_158 = 6'h1d == L0Index ? io_FromL1 : L0Memory_29; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_159 = 6'h1e == L0Index ? io_FromL1 : L0Memory_30; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_160 = 6'h1f == L0Index ? io_FromL1 : L0Memory_31; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_161 = 6'h20 == L0Index ? io_FromL1 : L0Memory_32; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_162 = 6'h21 == L0Index ? io_FromL1 : L0Memory_33; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_163 = 6'h22 == L0Index ? io_FromL1 : L0Memory_34; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_164 = 6'h23 == L0Index ? io_FromL1 : L0Memory_35; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_165 = 6'h24 == L0Index ? io_FromL1 : L0Memory_36; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_166 = 6'h25 == L0Index ? io_FromL1 : L0Memory_37; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_167 = 6'h26 == L0Index ? io_FromL1 : L0Memory_38; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_168 = 6'h27 == L0Index ? io_FromL1 : L0Memory_39; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_169 = 6'h28 == L0Index ? io_FromL1 : L0Memory_40; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_170 = 6'h29 == L0Index ? io_FromL1 : L0Memory_41; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_171 = 6'h2a == L0Index ? io_FromL1 : L0Memory_42; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_172 = 6'h2b == L0Index ? io_FromL1 : L0Memory_43; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_173 = 6'h2c == L0Index ? io_FromL1 : L0Memory_44; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_174 = 6'h2d == L0Index ? io_FromL1 : L0Memory_45; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_175 = 6'h2e == L0Index ? io_FromL1 : L0Memory_46; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_176 = 6'h2f == L0Index ? io_FromL1 : L0Memory_47; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_177 = 6'h30 == L0Index ? io_FromL1 : L0Memory_48; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_178 = 6'h31 == L0Index ? io_FromL1 : L0Memory_49; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_179 = 6'h32 == L0Index ? io_FromL1 : L0Memory_50; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_180 = 6'h33 == L0Index ? io_FromL1 : L0Memory_51; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_181 = 6'h34 == L0Index ? io_FromL1 : L0Memory_52; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_182 = 6'h35 == L0Index ? io_FromL1 : L0Memory_53; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_183 = 6'h36 == L0Index ? io_FromL1 : L0Memory_54; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_184 = 6'h37 == L0Index ? io_FromL1 : L0Memory_55; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_185 = 6'h38 == L0Index ? io_FromL1 : L0Memory_56; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_186 = 6'h39 == L0Index ? io_FromL1 : L0Memory_57; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_187 = 6'h3a == L0Index ? io_FromL1 : L0Memory_58; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_188 = 6'h3b == L0Index ? io_FromL1 : L0Memory_59; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_189 = 6'h3c == L0Index ? io_FromL1 : L0Memory_60; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_190 = 6'h3d == L0Index ? io_FromL1 : L0Memory_61; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_191 = 6'h3e == L0Index ? io_FromL1 : L0Memory_62; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_192 = 6'h3f == L0Index ? io_FromL1 : L0Memory_63; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_193 = 7'h40 == _GEN_793 ? io_FromL1 : L0Memory_64; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_194 = 7'h41 == _GEN_793 ? io_FromL1 : L0Memory_65; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_195 = 7'h42 == _GEN_793 ? io_FromL1 : L0Memory_66; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_196 = 7'h43 == _GEN_793 ? io_FromL1 : L0Memory_67; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_197 = 7'h44 == _GEN_793 ? io_FromL1 : L0Memory_68; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_198 = 7'h45 == _GEN_793 ? io_FromL1 : L0Memory_69; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_199 = 7'h46 == _GEN_793 ? io_FromL1 : L0Memory_70; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_200 = 7'h47 == _GEN_793 ? io_FromL1 : L0Memory_71; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_201 = 7'h48 == _GEN_793 ? io_FromL1 : L0Memory_72; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_202 = 7'h49 == _GEN_793 ? io_FromL1 : L0Memory_73; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_203 = 7'h4a == _GEN_793 ? io_FromL1 : L0Memory_74; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_204 = 7'h4b == _GEN_793 ? io_FromL1 : L0Memory_75; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_205 = 7'h4c == _GEN_793 ? io_FromL1 : L0Memory_76; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_206 = 7'h4d == _GEN_793 ? io_FromL1 : L0Memory_77; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_207 = 7'h4e == _GEN_793 ? io_FromL1 : L0Memory_78; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_208 = 7'h4f == _GEN_793 ? io_FromL1 : L0Memory_79; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_209 = 7'h50 == _GEN_793 ? io_FromL1 : L0Memory_80; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_210 = 7'h51 == _GEN_793 ? io_FromL1 : L0Memory_81; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_211 = 7'h52 == _GEN_793 ? io_FromL1 : L0Memory_82; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_212 = 7'h53 == _GEN_793 ? io_FromL1 : L0Memory_83; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_213 = 7'h54 == _GEN_793 ? io_FromL1 : L0Memory_84; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_214 = 7'h55 == _GEN_793 ? io_FromL1 : L0Memory_85; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_215 = 7'h56 == _GEN_793 ? io_FromL1 : L0Memory_86; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_216 = 7'h57 == _GEN_793 ? io_FromL1 : L0Memory_87; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_217 = 7'h58 == _GEN_793 ? io_FromL1 : L0Memory_88; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_218 = 7'h59 == _GEN_793 ? io_FromL1 : L0Memory_89; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_219 = 7'h5a == _GEN_793 ? io_FromL1 : L0Memory_90; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_220 = 7'h5b == _GEN_793 ? io_FromL1 : L0Memory_91; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_221 = 7'h5c == _GEN_793 ? io_FromL1 : L0Memory_92; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_222 = 7'h5d == _GEN_793 ? io_FromL1 : L0Memory_93; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_223 = 7'h5e == _GEN_793 ? io_FromL1 : L0Memory_94; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_224 = 7'h5f == _GEN_793 ? io_FromL1 : L0Memory_95; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_225 = 7'h60 == _GEN_793 ? io_FromL1 : L0Memory_96; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_226 = 7'h61 == _GEN_793 ? io_FromL1 : L0Memory_97; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_227 = 7'h62 == _GEN_793 ? io_FromL1 : L0Memory_98; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_228 = 7'h63 == _GEN_793 ? io_FromL1 : L0Memory_99; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [5:0] _L0Index_T_2 = L0Index + 6'h1; // @[PEArray.scala 200:28]
  wire [15:0] _GEN_229 = count >= 10'h1 & count <= _T_27 ? _GEN_129 : L0Memory_0; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_230 = count >= 10'h1 & count <= _T_27 ? _GEN_130 : L0Memory_1; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_231 = count >= 10'h1 & count <= _T_27 ? _GEN_131 : L0Memory_2; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_232 = count >= 10'h1 & count <= _T_27 ? _GEN_132 : L0Memory_3; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_233 = count >= 10'h1 & count <= _T_27 ? _GEN_133 : L0Memory_4; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_234 = count >= 10'h1 & count <= _T_27 ? _GEN_134 : L0Memory_5; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_235 = count >= 10'h1 & count <= _T_27 ? _GEN_135 : L0Memory_6; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_236 = count >= 10'h1 & count <= _T_27 ? _GEN_136 : L0Memory_7; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_237 = count >= 10'h1 & count <= _T_27 ? _GEN_137 : L0Memory_8; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_238 = count >= 10'h1 & count <= _T_27 ? _GEN_138 : L0Memory_9; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_239 = count >= 10'h1 & count <= _T_27 ? _GEN_139 : L0Memory_10; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_240 = count >= 10'h1 & count <= _T_27 ? _GEN_140 : L0Memory_11; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_241 = count >= 10'h1 & count <= _T_27 ? _GEN_141 : L0Memory_12; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_242 = count >= 10'h1 & count <= _T_27 ? _GEN_142 : L0Memory_13; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_243 = count >= 10'h1 & count <= _T_27 ? _GEN_143 : L0Memory_14; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_244 = count >= 10'h1 & count <= _T_27 ? _GEN_144 : L0Memory_15; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_245 = count >= 10'h1 & count <= _T_27 ? _GEN_145 : L0Memory_16; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_246 = count >= 10'h1 & count <= _T_27 ? _GEN_146 : L0Memory_17; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_247 = count >= 10'h1 & count <= _T_27 ? _GEN_147 : L0Memory_18; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_248 = count >= 10'h1 & count <= _T_27 ? _GEN_148 : L0Memory_19; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_249 = count >= 10'h1 & count <= _T_27 ? _GEN_149 : L0Memory_20; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_250 = count >= 10'h1 & count <= _T_27 ? _GEN_150 : L0Memory_21; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_251 = count >= 10'h1 & count <= _T_27 ? _GEN_151 : L0Memory_22; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_252 = count >= 10'h1 & count <= _T_27 ? _GEN_152 : L0Memory_23; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_253 = count >= 10'h1 & count <= _T_27 ? _GEN_153 : L0Memory_24; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_254 = count >= 10'h1 & count <= _T_27 ? _GEN_154 : L0Memory_25; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_255 = count >= 10'h1 & count <= _T_27 ? _GEN_155 : L0Memory_26; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_256 = count >= 10'h1 & count <= _T_27 ? _GEN_156 : L0Memory_27; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_257 = count >= 10'h1 & count <= _T_27 ? _GEN_157 : L0Memory_28; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_258 = count >= 10'h1 & count <= _T_27 ? _GEN_158 : L0Memory_29; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_259 = count >= 10'h1 & count <= _T_27 ? _GEN_159 : L0Memory_30; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_260 = count >= 10'h1 & count <= _T_27 ? _GEN_160 : L0Memory_31; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_261 = count >= 10'h1 & count <= _T_27 ? _GEN_161 : L0Memory_32; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_262 = count >= 10'h1 & count <= _T_27 ? _GEN_162 : L0Memory_33; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_263 = count >= 10'h1 & count <= _T_27 ? _GEN_163 : L0Memory_34; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_264 = count >= 10'h1 & count <= _T_27 ? _GEN_164 : L0Memory_35; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_265 = count >= 10'h1 & count <= _T_27 ? _GEN_165 : L0Memory_36; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_266 = count >= 10'h1 & count <= _T_27 ? _GEN_166 : L0Memory_37; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_267 = count >= 10'h1 & count <= _T_27 ? _GEN_167 : L0Memory_38; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_268 = count >= 10'h1 & count <= _T_27 ? _GEN_168 : L0Memory_39; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_269 = count >= 10'h1 & count <= _T_27 ? _GEN_169 : L0Memory_40; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_270 = count >= 10'h1 & count <= _T_27 ? _GEN_170 : L0Memory_41; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_271 = count >= 10'h1 & count <= _T_27 ? _GEN_171 : L0Memory_42; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_272 = count >= 10'h1 & count <= _T_27 ? _GEN_172 : L0Memory_43; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_273 = count >= 10'h1 & count <= _T_27 ? _GEN_173 : L0Memory_44; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_274 = count >= 10'h1 & count <= _T_27 ? _GEN_174 : L0Memory_45; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_275 = count >= 10'h1 & count <= _T_27 ? _GEN_175 : L0Memory_46; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_276 = count >= 10'h1 & count <= _T_27 ? _GEN_176 : L0Memory_47; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_277 = count >= 10'h1 & count <= _T_27 ? _GEN_177 : L0Memory_48; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_278 = count >= 10'h1 & count <= _T_27 ? _GEN_178 : L0Memory_49; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_279 = count >= 10'h1 & count <= _T_27 ? _GEN_179 : L0Memory_50; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_280 = count >= 10'h1 & count <= _T_27 ? _GEN_180 : L0Memory_51; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_281 = count >= 10'h1 & count <= _T_27 ? _GEN_181 : L0Memory_52; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_282 = count >= 10'h1 & count <= _T_27 ? _GEN_182 : L0Memory_53; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_283 = count >= 10'h1 & count <= _T_27 ? _GEN_183 : L0Memory_54; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_284 = count >= 10'h1 & count <= _T_27 ? _GEN_184 : L0Memory_55; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_285 = count >= 10'h1 & count <= _T_27 ? _GEN_185 : L0Memory_56; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_286 = count >= 10'h1 & count <= _T_27 ? _GEN_186 : L0Memory_57; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_287 = count >= 10'h1 & count <= _T_27 ? _GEN_187 : L0Memory_58; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_288 = count >= 10'h1 & count <= _T_27 ? _GEN_188 : L0Memory_59; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_289 = count >= 10'h1 & count <= _T_27 ? _GEN_189 : L0Memory_60; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_290 = count >= 10'h1 & count <= _T_27 ? _GEN_190 : L0Memory_61; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_291 = count >= 10'h1 & count <= _T_27 ? _GEN_191 : L0Memory_62; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_292 = count >= 10'h1 & count <= _T_27 ? _GEN_192 : L0Memory_63; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_293 = count >= 10'h1 & count <= _T_27 ? _GEN_193 : L0Memory_64; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_294 = count >= 10'h1 & count <= _T_27 ? _GEN_194 : L0Memory_65; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_295 = count >= 10'h1 & count <= _T_27 ? _GEN_195 : L0Memory_66; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_296 = count >= 10'h1 & count <= _T_27 ? _GEN_196 : L0Memory_67; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_297 = count >= 10'h1 & count <= _T_27 ? _GEN_197 : L0Memory_68; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_298 = count >= 10'h1 & count <= _T_27 ? _GEN_198 : L0Memory_69; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_299 = count >= 10'h1 & count <= _T_27 ? _GEN_199 : L0Memory_70; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_300 = count >= 10'h1 & count <= _T_27 ? _GEN_200 : L0Memory_71; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_301 = count >= 10'h1 & count <= _T_27 ? _GEN_201 : L0Memory_72; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_302 = count >= 10'h1 & count <= _T_27 ? _GEN_202 : L0Memory_73; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_303 = count >= 10'h1 & count <= _T_27 ? _GEN_203 : L0Memory_74; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_304 = count >= 10'h1 & count <= _T_27 ? _GEN_204 : L0Memory_75; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_305 = count >= 10'h1 & count <= _T_27 ? _GEN_205 : L0Memory_76; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_306 = count >= 10'h1 & count <= _T_27 ? _GEN_206 : L0Memory_77; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_307 = count >= 10'h1 & count <= _T_27 ? _GEN_207 : L0Memory_78; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_308 = count >= 10'h1 & count <= _T_27 ? _GEN_208 : L0Memory_79; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_309 = count >= 10'h1 & count <= _T_27 ? _GEN_209 : L0Memory_80; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_310 = count >= 10'h1 & count <= _T_27 ? _GEN_210 : L0Memory_81; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_311 = count >= 10'h1 & count <= _T_27 ? _GEN_211 : L0Memory_82; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_312 = count >= 10'h1 & count <= _T_27 ? _GEN_212 : L0Memory_83; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_313 = count >= 10'h1 & count <= _T_27 ? _GEN_213 : L0Memory_84; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_314 = count >= 10'h1 & count <= _T_27 ? _GEN_214 : L0Memory_85; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_315 = count >= 10'h1 & count <= _T_27 ? _GEN_215 : L0Memory_86; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_316 = count >= 10'h1 & count <= _T_27 ? _GEN_216 : L0Memory_87; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_317 = count >= 10'h1 & count <= _T_27 ? _GEN_217 : L0Memory_88; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_318 = count >= 10'h1 & count <= _T_27 ? _GEN_218 : L0Memory_89; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_319 = count >= 10'h1 & count <= _T_27 ? _GEN_219 : L0Memory_90; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_320 = count >= 10'h1 & count <= _T_27 ? _GEN_220 : L0Memory_91; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_321 = count >= 10'h1 & count <= _T_27 ? _GEN_221 : L0Memory_92; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_322 = count >= 10'h1 & count <= _T_27 ? _GEN_222 : L0Memory_93; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_323 = count >= 10'h1 & count <= _T_27 ? _GEN_223 : L0Memory_94; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_324 = count >= 10'h1 & count <= _T_27 ? _GEN_224 : L0Memory_95; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_325 = count >= 10'h1 & count <= _T_27 ? _GEN_225 : L0Memory_96; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_326 = count >= 10'h1 & count <= _T_27 ? _GEN_226 : L0Memory_97; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_327 = count >= 10'h1 & count <= _T_27 ? _GEN_227 : L0Memory_98; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_328 = count >= 10'h1 & count <= _T_27 ? _GEN_228 : L0Memory_99; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [5:0] _GEN_329 = count >= 10'h1 & count <= _T_27 ? _L0Index_T_2 : _GEN_128; // @[PEArray.scala 198:59 PEArray.scala 200:17]
  wire [9:0] _GEN_330 = _T_24 ? 10'h0 : _GEN_127; // @[PEArray.scala 202:32 PEArray.scala 203:15]
  wire [2:0] _GEN_331 = _T_24 ? 3'h0 : state; // @[PEArray.scala 202:32 PEArray.scala 204:15 PEArray.scala 100:22]
  wire [9:0] _GEN_865 = {{4'd0}, GRU_out_width}; // @[PEArray.scala 220:19]
  wire [9:0] _GEN_0 = count % _GEN_865; // @[PEArray.scala 220:19]
  wire [5:0] _T_36 = _GEN_0[5:0]; // @[PEArray.scala 220:19]
  wire [5:0] _T_38 = GRU_out_width - 6'h1; // @[PEArray.scala 220:55]
  wire [5:0] _GEN_334 = _T_36 == _T_38 ? _L0Index_T_2 : 6'h0; // @[PEArray.scala 220:62 PEArray.scala 221:17 PEArray.scala 214:15]
  wire [5:0] _GEN_346 = _T_41 ? _GEN_334 : L0Index; // @[Conditional.scala 39:67 PEArray.scala 39:24]
  wire [9:0] _GEN_347 = _T_41 ? _GEN_330 : count; // @[Conditional.scala 39:67 PEArray.scala 101:22]
  wire [2:0] _GEN_348 = _T_41 ? _GEN_331 : state; // @[Conditional.scala 39:67 PEArray.scala 100:22]
  wire [5:0] _GEN_353 = _T_31 ? _GEN_334 : _GEN_346; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_354 = _T_31 ? _GEN_330 : _GEN_347; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_355 = _T_31 ? _GEN_331 : _GEN_348; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_356 = _T_22 ? _GEN_330 : _GEN_354; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_357 = _T_22 ? _GEN_329 : _GEN_353; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_458 = _T_22 ? _GEN_331 : _GEN_355; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_690 = _T_3 ? _GEN_118 : {{2'd0}, GRU_out_width}; // @[Conditional.scala 40:58 PEArray.scala 104:26]
  FP16MulAdder FP16MAC ( // @[PEArray.scala 72:23]
    .io_a(FP16MAC_io_a),
    .io_b(FP16MAC_io_b),
    .io_c(FP16MAC_io_c),
    .io_out(FP16MAC_io_out)
  );
  assign io_ToRightPE = mux3out_reg; // @[PEArray.scala 95:16]
  assign io_ToBelowPE = mux2out_reg; // @[PEArray.scala 94:16]
  assign FP16MAC_io_a = sel1 ? io_FromL1 : io_FromLeftPE; // @[PEArray.scala 50:14 PEArray.scala 50:23 PEArray.scala 51:24]
  assign FP16MAC_io_b = sel5 ? mux4out : _GEN_105; // @[PEArray.scala 77:13 PEArray.scala 78:18 PEArray.scala 81:18]
  assign FP16MAC_io_c = sel5 ? _GEN_105 : mux4out; // @[PEArray.scala 77:13 PEArray.scala 79:18 PEArray.scala 82:18]
  always @(posedge clock) begin
    if (reset) begin // @[PEArray.scala 39:24]
      L0Index <= 6'h0; // @[PEArray.scala 39:24]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h0; // @[PEArray.scala 159:15]
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        L0Index <= 6'hb; // @[PEArray.scala 181:15]
      end else begin
        L0Index <= _GEN_357;
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_0 <= _GEN_229;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_1 <= _GEN_230;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_2 <= _GEN_231;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_3 <= _GEN_232;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_4 <= _GEN_233;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_5 <= _GEN_234;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_6 <= _GEN_235;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_7 <= _GEN_236;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_8 <= _GEN_237;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_9 <= _GEN_238;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_10 <= _GEN_239;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_11 <= _GEN_240;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_12 <= _GEN_241;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_13 <= _GEN_242;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_14 <= _GEN_243;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_15 <= _GEN_244;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_16 <= _GEN_245;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_17 <= _GEN_246;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_18 <= _GEN_247;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_19 <= _GEN_248;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_20 <= _GEN_249;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_21 <= _GEN_250;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_22 <= _GEN_251;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_23 <= _GEN_252;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_24 <= _GEN_253;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_25 <= _GEN_254;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_26 <= _GEN_255;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_27 <= _GEN_256;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_28 <= _GEN_257;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_29 <= _GEN_258;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_30 <= _GEN_259;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_31 <= _GEN_260;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_32 <= _GEN_261;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_33 <= _GEN_262;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_34 <= _GEN_263;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_35 <= _GEN_264;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_36 <= _GEN_265;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_37 <= _GEN_266;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_38 <= _GEN_267;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_39 <= _GEN_268;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_40 <= _GEN_269;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_41 <= _GEN_270;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_42 <= _GEN_271;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_43 <= _GEN_272;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_44 <= _GEN_273;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_45 <= _GEN_274;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_46 <= _GEN_275;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_47 <= _GEN_276;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_48 <= _GEN_277;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_49 <= _GEN_278;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_50 <= _GEN_279;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_51 <= _GEN_280;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_52 <= _GEN_281;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_53 <= _GEN_282;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_54 <= _GEN_283;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_55 <= _GEN_284;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_56 <= _GEN_285;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_57 <= _GEN_286;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_58 <= _GEN_287;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_59 <= _GEN_288;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_60 <= _GEN_289;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_61 <= _GEN_290;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_62 <= _GEN_291;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_63 <= _GEN_292;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_64 <= _GEN_293;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_65 <= _GEN_294;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_66 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_67 <= _GEN_296;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_68 <= _GEN_297;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_69 <= _GEN_298;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_70 <= _GEN_299;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_71 <= _GEN_300;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_72 <= _GEN_301;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_73 <= _GEN_302;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_74 <= _GEN_303;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_75 <= _GEN_304;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_76 <= _GEN_305;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_77 <= _GEN_306;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_78 <= _GEN_307;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_79 <= _GEN_308;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_80 <= _GEN_309;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_81 <= _GEN_310;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_82 <= _GEN_311;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_83 <= _GEN_312;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_84 <= _GEN_313;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_85 <= _GEN_314;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_86 <= _GEN_315;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_87 <= _GEN_316;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_88 <= _GEN_317;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_89 <= _GEN_318;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_90 <= _GEN_319;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_91 <= _GEN_320;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_92 <= _GEN_321;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_93 <= _GEN_322;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_94 <= _GEN_323;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_95 <= _GEN_324;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_96 <= _GEN_325;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_97 <= _GEN_326;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_98 <= _GEN_327;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_99 <= _GEN_328;
          end
        end
      end
    end
    if (reset) begin // @[PEArray.scala 100:22]
      state <= 3'h0; // @[PEArray.scala 100:22]
    end else if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[3]) begin // @[PEArray.scala 116:57]
        state <= 3'h1;
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      if (count == 10'h33) begin // @[PEArray.scala 164:27]
        state <= 3'h0; // @[PEArray.scala 166:15]
      end
    end else if (_T_16) begin // @[Conditional.scala 39:67]
      state <= _GEN_126;
    end else begin
      state <= _GEN_458;
    end
    if (reset) begin // @[PEArray.scala 90:28]
      mux2out_reg <= 16'h0; // @[PEArray.scala 90:28]
    end else begin
      mux2out_reg <= MAC_out; // @[PEArray.scala 90:28]
    end
    if (reset) begin // @[PEArray.scala 91:28]
      mux3out_reg <= 16'h0; // @[PEArray.scala 91:28]
    end else if (sel3) begin // @[PEArray.scala 56:14]
      mux3out_reg <= MAC_out; // @[PEArray.scala 56:23]
    end else if (sel1) begin // @[PEArray.scala 50:14]
      mux3out_reg <= io_FromL1; // @[PEArray.scala 50:23]
    end else begin
      mux3out_reg <= io_FromLeftPE; // @[PEArray.scala 51:24]
    end
    if (reset) begin // @[PEArray.scala 101:22]
      count <= 10'h0; // @[PEArray.scala 101:22]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        if (count == 10'h33) begin // @[PEArray.scala 164:27]
          count <= 10'h0; // @[PEArray.scala 165:15]
        end else begin
          count <= _GEN_120;
        end
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        count <= _GEN_125;
      end else begin
        count <= _GEN_356;
      end
    end
    GRU_out_width <= _GEN_690[5:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  L0Index = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  L0Memory_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  L0Memory_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  L0Memory_2 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  L0Memory_3 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  L0Memory_4 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  L0Memory_5 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  L0Memory_6 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  L0Memory_7 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  L0Memory_8 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  L0Memory_9 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  L0Memory_10 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  L0Memory_11 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  L0Memory_12 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  L0Memory_13 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  L0Memory_14 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  L0Memory_15 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  L0Memory_16 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  L0Memory_17 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  L0Memory_18 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  L0Memory_19 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  L0Memory_20 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  L0Memory_21 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  L0Memory_22 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  L0Memory_23 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  L0Memory_24 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  L0Memory_25 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  L0Memory_26 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  L0Memory_27 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  L0Memory_28 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  L0Memory_29 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  L0Memory_30 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  L0Memory_31 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  L0Memory_32 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  L0Memory_33 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  L0Memory_34 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  L0Memory_35 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  L0Memory_36 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  L0Memory_37 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  L0Memory_38 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  L0Memory_39 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  L0Memory_40 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  L0Memory_41 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  L0Memory_42 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  L0Memory_43 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  L0Memory_44 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  L0Memory_45 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  L0Memory_46 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  L0Memory_47 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  L0Memory_48 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  L0Memory_49 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  L0Memory_50 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  L0Memory_51 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  L0Memory_52 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  L0Memory_53 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  L0Memory_54 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  L0Memory_55 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  L0Memory_56 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  L0Memory_57 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  L0Memory_58 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  L0Memory_59 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  L0Memory_60 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  L0Memory_61 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  L0Memory_62 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  L0Memory_63 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  L0Memory_64 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  L0Memory_65 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  L0Memory_66 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  L0Memory_67 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  L0Memory_68 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  L0Memory_69 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  L0Memory_70 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  L0Memory_71 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  L0Memory_72 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  L0Memory_73 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  L0Memory_74 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  L0Memory_75 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  L0Memory_76 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  L0Memory_77 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  L0Memory_78 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  L0Memory_79 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  L0Memory_80 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  L0Memory_81 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  L0Memory_82 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  L0Memory_83 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  L0Memory_84 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  L0Memory_85 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  L0Memory_86 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  L0Memory_87 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  L0Memory_88 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  L0Memory_89 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  L0Memory_90 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  L0Memory_91 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  L0Memory_92 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  L0Memory_93 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  L0Memory_94 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  L0Memory_95 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  L0Memory_96 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  L0Memory_97 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  L0Memory_98 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  L0Memory_99 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  state = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  mux2out_reg = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  mux3out_reg = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  count = _RAND_104[9:0];
  _RAND_105 = {1{`RANDOM}};
  GRU_out_width = _RAND_105[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PE_25(
  input         clock,
  input         reset,
  input  [15:0] io_FromAbovePE,
  input  [15:0] io_FromLeftPE,
  input  [15:0] io_FromL1,
  input  [11:0] io_control_signal_mask,
  output [15:0] io_ToRightPE,
  output [15:0] io_ToBelowPE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] FP16MAC_io_a; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_b; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_c; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_out; // @[PEArray.scala 72:23]
  reg [5:0] L0Index; // @[PEArray.scala 39:24]
  reg [15:0] L0Memory_0; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_1; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_2; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_3; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_4; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_5; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_6; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_7; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_8; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_9; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_10; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_11; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_12; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_13; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_14; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_15; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_16; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_17; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_18; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_19; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_20; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_21; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_22; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_23; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_24; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_25; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_26; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_27; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_28; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_29; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_30; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_31; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_32; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_33; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_34; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_35; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_36; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_37; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_38; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_39; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_40; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_41; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_42; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_43; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_44; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_45; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_46; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_47; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_48; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_49; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_50; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_51; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_52; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_53; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_54; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_55; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_56; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_57; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_58; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_59; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_60; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_61; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_62; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_63; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_64; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_65; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_66; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_67; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_68; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_69; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_70; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_71; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_72; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_73; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_74; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_75; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_76; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_77; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_78; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_79; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_80; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_81; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_82; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_83; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_84; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_85; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_86; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_87; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_88; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_89; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_90; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_91; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_92; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_93; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_94; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_95; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_96; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_97; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_98; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_99; // @[PEArray.scala 40:21]
  reg [2:0] state; // @[PEArray.scala 100:22]
  wire  _T_3 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_12 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_16 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_22 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_31 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_41 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_342 = _T_41 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 231:12 PEArray.scala 32:8]
  wire  _GEN_349 = _T_31 ? 1'h0 : _GEN_342; // @[Conditional.scala 39:67 PEArray.scala 208:12]
  wire  _GEN_459 = _T_22 | _GEN_349; // @[Conditional.scala 39:67 PEArray.scala 32:8]
  wire  _GEN_463 = _T_16 ? 1'h0 : _GEN_459; // @[Conditional.scala 39:67]
  wire  _GEN_572 = _T_12 | _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 149:12]
  wire  sel1 = _T_3 | _GEN_572; // @[Conditional.scala 40:58 PEArray.scala 108:12]
  wire [15:0] MAC_out = FP16MAC_io_out; // @[PEArray.scala 47:21 PEArray.scala 85:11]
  wire  _GEN_465 = _T_16 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 177:12]
  wire  _GEN_580 = _T_12 | _GEN_465; // @[Conditional.scala 39:67 PEArray.scala 34:8]
  wire  sel3 = _T_3 | _GEN_580; // @[Conditional.scala 40:58 PEArray.scala 110:12]
  wire [1:0] _GEN_344 = _T_41 ? 2'h2 : 2'h0; // @[Conditional.scala 39:67 PEArray.scala 233:12 PEArray.scala 35:8]
  wire [1:0] _GEN_351 = _T_31 ? 2'h2 : _GEN_344; // @[Conditional.scala 39:67 PEArray.scala 210:12]
  wire [1:0] _GEN_461 = _T_22 ? 2'h0 : _GEN_351; // @[Conditional.scala 39:67 PEArray.scala 35:8]
  wire [1:0] _GEN_466 = _T_16 ? 2'h0 : _GEN_461; // @[Conditional.scala 39:67 PEArray.scala 178:12]
  wire [1:0] _GEN_574 = _T_12 ? 2'h1 : _GEN_466; // @[Conditional.scala 39:67]
  wire [1:0] sel4 = _T_3 ? 2'h0 : _GEN_574; // @[Conditional.scala 40:58 PEArray.scala 111:12]
  wire [15:0] _GEN_3 = sel4 == 2'h2 ? io_FromL1 : 16'h0; // @[PEArray.scala 65:28 PEArray.scala 66:15 PEArray.scala 69:15]
  wire [15:0] _GEN_4 = sel4 == 2'h1 ? io_FromAbovePE : _GEN_3; // @[PEArray.scala 62:28 PEArray.scala 63:15]
  wire [15:0] mux4out = sel4 == 2'h0 ? 16'h0 : _GEN_4; // @[PEArray.scala 59:22 PEArray.scala 60:13]
  wire [15:0] _GEN_7 = 6'h1 == L0Index ? L0Memory_1 : L0Memory_0; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_8 = 6'h2 == L0Index ? L0Memory_2 : _GEN_7; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_9 = 6'h3 == L0Index ? L0Memory_3 : _GEN_8; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_10 = 6'h4 == L0Index ? L0Memory_4 : _GEN_9; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_11 = 6'h5 == L0Index ? L0Memory_5 : _GEN_10; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_12 = 6'h6 == L0Index ? L0Memory_6 : _GEN_11; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_13 = 6'h7 == L0Index ? L0Memory_7 : _GEN_12; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_14 = 6'h8 == L0Index ? L0Memory_8 : _GEN_13; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_15 = 6'h9 == L0Index ? L0Memory_9 : _GEN_14; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_16 = 6'ha == L0Index ? L0Memory_10 : _GEN_15; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_17 = 6'hb == L0Index ? L0Memory_11 : _GEN_16; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_18 = 6'hc == L0Index ? L0Memory_12 : _GEN_17; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_19 = 6'hd == L0Index ? L0Memory_13 : _GEN_18; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_20 = 6'he == L0Index ? L0Memory_14 : _GEN_19; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_21 = 6'hf == L0Index ? L0Memory_15 : _GEN_20; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_22 = 6'h10 == L0Index ? L0Memory_16 : _GEN_21; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_23 = 6'h11 == L0Index ? L0Memory_17 : _GEN_22; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_24 = 6'h12 == L0Index ? L0Memory_18 : _GEN_23; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_25 = 6'h13 == L0Index ? L0Memory_19 : _GEN_24; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_26 = 6'h14 == L0Index ? L0Memory_20 : _GEN_25; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_27 = 6'h15 == L0Index ? L0Memory_21 : _GEN_26; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_28 = 6'h16 == L0Index ? L0Memory_22 : _GEN_27; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_29 = 6'h17 == L0Index ? L0Memory_23 : _GEN_28; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_30 = 6'h18 == L0Index ? L0Memory_24 : _GEN_29; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_31 = 6'h19 == L0Index ? L0Memory_25 : _GEN_30; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_32 = 6'h1a == L0Index ? L0Memory_26 : _GEN_31; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_33 = 6'h1b == L0Index ? L0Memory_27 : _GEN_32; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_34 = 6'h1c == L0Index ? L0Memory_28 : _GEN_33; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_35 = 6'h1d == L0Index ? L0Memory_29 : _GEN_34; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_36 = 6'h1e == L0Index ? L0Memory_30 : _GEN_35; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_37 = 6'h1f == L0Index ? L0Memory_31 : _GEN_36; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_38 = 6'h20 == L0Index ? L0Memory_32 : _GEN_37; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_39 = 6'h21 == L0Index ? L0Memory_33 : _GEN_38; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_40 = 6'h22 == L0Index ? L0Memory_34 : _GEN_39; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_41 = 6'h23 == L0Index ? L0Memory_35 : _GEN_40; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_42 = 6'h24 == L0Index ? L0Memory_36 : _GEN_41; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_43 = 6'h25 == L0Index ? L0Memory_37 : _GEN_42; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_44 = 6'h26 == L0Index ? L0Memory_38 : _GEN_43; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_45 = 6'h27 == L0Index ? L0Memory_39 : _GEN_44; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_46 = 6'h28 == L0Index ? L0Memory_40 : _GEN_45; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_47 = 6'h29 == L0Index ? L0Memory_41 : _GEN_46; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_48 = 6'h2a == L0Index ? L0Memory_42 : _GEN_47; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_49 = 6'h2b == L0Index ? L0Memory_43 : _GEN_48; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_50 = 6'h2c == L0Index ? L0Memory_44 : _GEN_49; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_51 = 6'h2d == L0Index ? L0Memory_45 : _GEN_50; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_52 = 6'h2e == L0Index ? L0Memory_46 : _GEN_51; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_53 = 6'h2f == L0Index ? L0Memory_47 : _GEN_52; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_54 = 6'h30 == L0Index ? L0Memory_48 : _GEN_53; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_55 = 6'h31 == L0Index ? L0Memory_49 : _GEN_54; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_56 = 6'h32 == L0Index ? L0Memory_50 : _GEN_55; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_57 = 6'h33 == L0Index ? L0Memory_51 : _GEN_56; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_58 = 6'h34 == L0Index ? L0Memory_52 : _GEN_57; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_59 = 6'h35 == L0Index ? L0Memory_53 : _GEN_58; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_60 = 6'h36 == L0Index ? L0Memory_54 : _GEN_59; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_61 = 6'h37 == L0Index ? L0Memory_55 : _GEN_60; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_62 = 6'h38 == L0Index ? L0Memory_56 : _GEN_61; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_63 = 6'h39 == L0Index ? L0Memory_57 : _GEN_62; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_64 = 6'h3a == L0Index ? L0Memory_58 : _GEN_63; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_65 = 6'h3b == L0Index ? L0Memory_59 : _GEN_64; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_66 = 6'h3c == L0Index ? L0Memory_60 : _GEN_65; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_67 = 6'h3d == L0Index ? L0Memory_61 : _GEN_66; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_68 = 6'h3e == L0Index ? L0Memory_62 : _GEN_67; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_69 = 6'h3f == L0Index ? L0Memory_63 : _GEN_68; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [6:0] _GEN_793 = {{1'd0}, L0Index}; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_70 = 7'h40 == _GEN_793 ? L0Memory_64 : _GEN_69; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_71 = 7'h41 == _GEN_793 ? L0Memory_65 : _GEN_70; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_72 = 7'h42 == _GEN_793 ? L0Memory_66 : _GEN_71; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_73 = 7'h43 == _GEN_793 ? L0Memory_67 : _GEN_72; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_74 = 7'h44 == _GEN_793 ? L0Memory_68 : _GEN_73; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_75 = 7'h45 == _GEN_793 ? L0Memory_69 : _GEN_74; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_76 = 7'h46 == _GEN_793 ? L0Memory_70 : _GEN_75; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_77 = 7'h47 == _GEN_793 ? L0Memory_71 : _GEN_76; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_78 = 7'h48 == _GEN_793 ? L0Memory_72 : _GEN_77; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_79 = 7'h49 == _GEN_793 ? L0Memory_73 : _GEN_78; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_80 = 7'h4a == _GEN_793 ? L0Memory_74 : _GEN_79; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_81 = 7'h4b == _GEN_793 ? L0Memory_75 : _GEN_80; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_82 = 7'h4c == _GEN_793 ? L0Memory_76 : _GEN_81; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_83 = 7'h4d == _GEN_793 ? L0Memory_77 : _GEN_82; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_84 = 7'h4e == _GEN_793 ? L0Memory_78 : _GEN_83; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_85 = 7'h4f == _GEN_793 ? L0Memory_79 : _GEN_84; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_86 = 7'h50 == _GEN_793 ? L0Memory_80 : _GEN_85; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_87 = 7'h51 == _GEN_793 ? L0Memory_81 : _GEN_86; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_88 = 7'h52 == _GEN_793 ? L0Memory_82 : _GEN_87; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_89 = 7'h53 == _GEN_793 ? L0Memory_83 : _GEN_88; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_90 = 7'h54 == _GEN_793 ? L0Memory_84 : _GEN_89; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_91 = 7'h55 == _GEN_793 ? L0Memory_85 : _GEN_90; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_92 = 7'h56 == _GEN_793 ? L0Memory_86 : _GEN_91; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_93 = 7'h57 == _GEN_793 ? L0Memory_87 : _GEN_92; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_94 = 7'h58 == _GEN_793 ? L0Memory_88 : _GEN_93; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_95 = 7'h59 == _GEN_793 ? L0Memory_89 : _GEN_94; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_96 = 7'h5a == _GEN_793 ? L0Memory_90 : _GEN_95; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_97 = 7'h5b == _GEN_793 ? L0Memory_91 : _GEN_96; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_98 = 7'h5c == _GEN_793 ? L0Memory_92 : _GEN_97; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_99 = 7'h5d == _GEN_793 ? L0Memory_93 : _GEN_98; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_100 = 7'h5e == _GEN_793 ? L0Memory_94 : _GEN_99; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_101 = 7'h5f == _GEN_793 ? L0Memory_95 : _GEN_100; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_102 = 7'h60 == _GEN_793 ? L0Memory_96 : _GEN_101; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_103 = 7'h61 == _GEN_793 ? L0Memory_97 : _GEN_102; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_104 = 7'h62 == _GEN_793 ? L0Memory_98 : _GEN_103; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_105 = 7'h63 == _GEN_793 ? L0Memory_99 : _GEN_104; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire  _GEN_575 = _T_12 ? 1'h0 : _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 157:12]
  wire  sel5 = _T_3 ? 1'h0 : _GEN_575; // @[Conditional.scala 40:58 PEArray.scala 112:12]
  reg [15:0] mux2out_reg; // @[PEArray.scala 90:28]
  reg [15:0] mux3out_reg; // @[PEArray.scala 91:28]
  reg [9:0] count; // @[PEArray.scala 101:22]
  reg [5:0] GRU_out_width; // @[PEArray.scala 104:26]
  wire [7:0] _GEN_118 = io_control_signal_mask[3] ? 8'h0 : {{2'd0}, GRU_out_width}; // @[PEArray.scala 116:57 PEArray.scala 145:23 PEArray.scala 104:26]
  wire [9:0] _count_T_1 = count + 10'h1; // @[PEArray.scala 162:24]
  wire [9:0] _GEN_120 = count != 10'h33 ? _count_T_1 : count; // @[PEArray.scala 161:27 PEArray.scala 162:15 PEArray.scala 101:22]
  wire [9:0] _GEN_124 = count != 10'h188 ? _count_T_1 : count; // @[PEArray.scala 183:28 PEArray.scala 184:15 PEArray.scala 101:22]
  wire [9:0] _GEN_125 = count == 10'h188 ? 10'h0 : _GEN_124; // @[PEArray.scala 186:28 PEArray.scala 187:15]
  wire [2:0] _GEN_126 = count == 10'h188 ? 3'h0 : state; // @[PEArray.scala 186:28 PEArray.scala 188:15 PEArray.scala 100:22]
  wire [9:0] _GEN_127 = count != 10'h0 ? _count_T_1 : count; // @[PEArray.scala 192:32 PEArray.scala 193:15 PEArray.scala 101:22]
  wire  _T_24 = count == 10'h0; // @[PEArray.scala 195:18]
  wire [5:0] _GEN_128 = count == 10'h0 ? 6'h0 : L0Index; // @[PEArray.scala 195:26 PEArray.scala 196:17 PEArray.scala 39:24]
  wire [9:0] _T_27 = 10'h0 - 10'h1; // @[PEArray.scala 198:51]
  wire [15:0] _GEN_129 = 6'h0 == L0Index ? io_FromL1 : L0Memory_0; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_130 = 6'h1 == L0Index ? io_FromL1 : L0Memory_1; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_131 = 6'h2 == L0Index ? io_FromL1 : L0Memory_2; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_132 = 6'h3 == L0Index ? io_FromL1 : L0Memory_3; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_133 = 6'h4 == L0Index ? io_FromL1 : L0Memory_4; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_134 = 6'h5 == L0Index ? io_FromL1 : L0Memory_5; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_135 = 6'h6 == L0Index ? io_FromL1 : L0Memory_6; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_136 = 6'h7 == L0Index ? io_FromL1 : L0Memory_7; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_137 = 6'h8 == L0Index ? io_FromL1 : L0Memory_8; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_138 = 6'h9 == L0Index ? io_FromL1 : L0Memory_9; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_139 = 6'ha == L0Index ? io_FromL1 : L0Memory_10; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_140 = 6'hb == L0Index ? io_FromL1 : L0Memory_11; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_141 = 6'hc == L0Index ? io_FromL1 : L0Memory_12; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_142 = 6'hd == L0Index ? io_FromL1 : L0Memory_13; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_143 = 6'he == L0Index ? io_FromL1 : L0Memory_14; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_144 = 6'hf == L0Index ? io_FromL1 : L0Memory_15; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_145 = 6'h10 == L0Index ? io_FromL1 : L0Memory_16; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_146 = 6'h11 == L0Index ? io_FromL1 : L0Memory_17; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_147 = 6'h12 == L0Index ? io_FromL1 : L0Memory_18; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_148 = 6'h13 == L0Index ? io_FromL1 : L0Memory_19; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_149 = 6'h14 == L0Index ? io_FromL1 : L0Memory_20; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_150 = 6'h15 == L0Index ? io_FromL1 : L0Memory_21; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_151 = 6'h16 == L0Index ? io_FromL1 : L0Memory_22; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_152 = 6'h17 == L0Index ? io_FromL1 : L0Memory_23; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_153 = 6'h18 == L0Index ? io_FromL1 : L0Memory_24; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_154 = 6'h19 == L0Index ? io_FromL1 : L0Memory_25; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_155 = 6'h1a == L0Index ? io_FromL1 : L0Memory_26; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_156 = 6'h1b == L0Index ? io_FromL1 : L0Memory_27; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_157 = 6'h1c == L0Index ? io_FromL1 : L0Memory_28; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_158 = 6'h1d == L0Index ? io_FromL1 : L0Memory_29; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_159 = 6'h1e == L0Index ? io_FromL1 : L0Memory_30; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_160 = 6'h1f == L0Index ? io_FromL1 : L0Memory_31; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_161 = 6'h20 == L0Index ? io_FromL1 : L0Memory_32; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_162 = 6'h21 == L0Index ? io_FromL1 : L0Memory_33; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_163 = 6'h22 == L0Index ? io_FromL1 : L0Memory_34; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_164 = 6'h23 == L0Index ? io_FromL1 : L0Memory_35; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_165 = 6'h24 == L0Index ? io_FromL1 : L0Memory_36; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_166 = 6'h25 == L0Index ? io_FromL1 : L0Memory_37; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_167 = 6'h26 == L0Index ? io_FromL1 : L0Memory_38; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_168 = 6'h27 == L0Index ? io_FromL1 : L0Memory_39; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_169 = 6'h28 == L0Index ? io_FromL1 : L0Memory_40; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_170 = 6'h29 == L0Index ? io_FromL1 : L0Memory_41; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_171 = 6'h2a == L0Index ? io_FromL1 : L0Memory_42; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_172 = 6'h2b == L0Index ? io_FromL1 : L0Memory_43; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_173 = 6'h2c == L0Index ? io_FromL1 : L0Memory_44; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_174 = 6'h2d == L0Index ? io_FromL1 : L0Memory_45; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_175 = 6'h2e == L0Index ? io_FromL1 : L0Memory_46; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_176 = 6'h2f == L0Index ? io_FromL1 : L0Memory_47; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_177 = 6'h30 == L0Index ? io_FromL1 : L0Memory_48; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_178 = 6'h31 == L0Index ? io_FromL1 : L0Memory_49; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_179 = 6'h32 == L0Index ? io_FromL1 : L0Memory_50; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_180 = 6'h33 == L0Index ? io_FromL1 : L0Memory_51; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_181 = 6'h34 == L0Index ? io_FromL1 : L0Memory_52; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_182 = 6'h35 == L0Index ? io_FromL1 : L0Memory_53; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_183 = 6'h36 == L0Index ? io_FromL1 : L0Memory_54; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_184 = 6'h37 == L0Index ? io_FromL1 : L0Memory_55; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_185 = 6'h38 == L0Index ? io_FromL1 : L0Memory_56; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_186 = 6'h39 == L0Index ? io_FromL1 : L0Memory_57; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_187 = 6'h3a == L0Index ? io_FromL1 : L0Memory_58; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_188 = 6'h3b == L0Index ? io_FromL1 : L0Memory_59; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_189 = 6'h3c == L0Index ? io_FromL1 : L0Memory_60; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_190 = 6'h3d == L0Index ? io_FromL1 : L0Memory_61; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_191 = 6'h3e == L0Index ? io_FromL1 : L0Memory_62; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_192 = 6'h3f == L0Index ? io_FromL1 : L0Memory_63; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_193 = 7'h40 == _GEN_793 ? io_FromL1 : L0Memory_64; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_194 = 7'h41 == _GEN_793 ? io_FromL1 : L0Memory_65; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_195 = 7'h42 == _GEN_793 ? io_FromL1 : L0Memory_66; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_196 = 7'h43 == _GEN_793 ? io_FromL1 : L0Memory_67; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_197 = 7'h44 == _GEN_793 ? io_FromL1 : L0Memory_68; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_198 = 7'h45 == _GEN_793 ? io_FromL1 : L0Memory_69; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_199 = 7'h46 == _GEN_793 ? io_FromL1 : L0Memory_70; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_200 = 7'h47 == _GEN_793 ? io_FromL1 : L0Memory_71; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_201 = 7'h48 == _GEN_793 ? io_FromL1 : L0Memory_72; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_202 = 7'h49 == _GEN_793 ? io_FromL1 : L0Memory_73; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_203 = 7'h4a == _GEN_793 ? io_FromL1 : L0Memory_74; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_204 = 7'h4b == _GEN_793 ? io_FromL1 : L0Memory_75; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_205 = 7'h4c == _GEN_793 ? io_FromL1 : L0Memory_76; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_206 = 7'h4d == _GEN_793 ? io_FromL1 : L0Memory_77; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_207 = 7'h4e == _GEN_793 ? io_FromL1 : L0Memory_78; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_208 = 7'h4f == _GEN_793 ? io_FromL1 : L0Memory_79; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_209 = 7'h50 == _GEN_793 ? io_FromL1 : L0Memory_80; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_210 = 7'h51 == _GEN_793 ? io_FromL1 : L0Memory_81; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_211 = 7'h52 == _GEN_793 ? io_FromL1 : L0Memory_82; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_212 = 7'h53 == _GEN_793 ? io_FromL1 : L0Memory_83; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_213 = 7'h54 == _GEN_793 ? io_FromL1 : L0Memory_84; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_214 = 7'h55 == _GEN_793 ? io_FromL1 : L0Memory_85; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_215 = 7'h56 == _GEN_793 ? io_FromL1 : L0Memory_86; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_216 = 7'h57 == _GEN_793 ? io_FromL1 : L0Memory_87; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_217 = 7'h58 == _GEN_793 ? io_FromL1 : L0Memory_88; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_218 = 7'h59 == _GEN_793 ? io_FromL1 : L0Memory_89; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_219 = 7'h5a == _GEN_793 ? io_FromL1 : L0Memory_90; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_220 = 7'h5b == _GEN_793 ? io_FromL1 : L0Memory_91; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_221 = 7'h5c == _GEN_793 ? io_FromL1 : L0Memory_92; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_222 = 7'h5d == _GEN_793 ? io_FromL1 : L0Memory_93; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_223 = 7'h5e == _GEN_793 ? io_FromL1 : L0Memory_94; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_224 = 7'h5f == _GEN_793 ? io_FromL1 : L0Memory_95; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_225 = 7'h60 == _GEN_793 ? io_FromL1 : L0Memory_96; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_226 = 7'h61 == _GEN_793 ? io_FromL1 : L0Memory_97; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_227 = 7'h62 == _GEN_793 ? io_FromL1 : L0Memory_98; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_228 = 7'h63 == _GEN_793 ? io_FromL1 : L0Memory_99; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [5:0] _L0Index_T_2 = L0Index + 6'h1; // @[PEArray.scala 200:28]
  wire [15:0] _GEN_229 = count >= 10'h1 & count <= _T_27 ? _GEN_129 : L0Memory_0; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_230 = count >= 10'h1 & count <= _T_27 ? _GEN_130 : L0Memory_1; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_231 = count >= 10'h1 & count <= _T_27 ? _GEN_131 : L0Memory_2; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_232 = count >= 10'h1 & count <= _T_27 ? _GEN_132 : L0Memory_3; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_233 = count >= 10'h1 & count <= _T_27 ? _GEN_133 : L0Memory_4; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_234 = count >= 10'h1 & count <= _T_27 ? _GEN_134 : L0Memory_5; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_235 = count >= 10'h1 & count <= _T_27 ? _GEN_135 : L0Memory_6; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_236 = count >= 10'h1 & count <= _T_27 ? _GEN_136 : L0Memory_7; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_237 = count >= 10'h1 & count <= _T_27 ? _GEN_137 : L0Memory_8; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_238 = count >= 10'h1 & count <= _T_27 ? _GEN_138 : L0Memory_9; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_239 = count >= 10'h1 & count <= _T_27 ? _GEN_139 : L0Memory_10; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_240 = count >= 10'h1 & count <= _T_27 ? _GEN_140 : L0Memory_11; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_241 = count >= 10'h1 & count <= _T_27 ? _GEN_141 : L0Memory_12; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_242 = count >= 10'h1 & count <= _T_27 ? _GEN_142 : L0Memory_13; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_243 = count >= 10'h1 & count <= _T_27 ? _GEN_143 : L0Memory_14; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_244 = count >= 10'h1 & count <= _T_27 ? _GEN_144 : L0Memory_15; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_245 = count >= 10'h1 & count <= _T_27 ? _GEN_145 : L0Memory_16; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_246 = count >= 10'h1 & count <= _T_27 ? _GEN_146 : L0Memory_17; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_247 = count >= 10'h1 & count <= _T_27 ? _GEN_147 : L0Memory_18; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_248 = count >= 10'h1 & count <= _T_27 ? _GEN_148 : L0Memory_19; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_249 = count >= 10'h1 & count <= _T_27 ? _GEN_149 : L0Memory_20; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_250 = count >= 10'h1 & count <= _T_27 ? _GEN_150 : L0Memory_21; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_251 = count >= 10'h1 & count <= _T_27 ? _GEN_151 : L0Memory_22; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_252 = count >= 10'h1 & count <= _T_27 ? _GEN_152 : L0Memory_23; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_253 = count >= 10'h1 & count <= _T_27 ? _GEN_153 : L0Memory_24; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_254 = count >= 10'h1 & count <= _T_27 ? _GEN_154 : L0Memory_25; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_255 = count >= 10'h1 & count <= _T_27 ? _GEN_155 : L0Memory_26; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_256 = count >= 10'h1 & count <= _T_27 ? _GEN_156 : L0Memory_27; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_257 = count >= 10'h1 & count <= _T_27 ? _GEN_157 : L0Memory_28; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_258 = count >= 10'h1 & count <= _T_27 ? _GEN_158 : L0Memory_29; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_259 = count >= 10'h1 & count <= _T_27 ? _GEN_159 : L0Memory_30; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_260 = count >= 10'h1 & count <= _T_27 ? _GEN_160 : L0Memory_31; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_261 = count >= 10'h1 & count <= _T_27 ? _GEN_161 : L0Memory_32; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_262 = count >= 10'h1 & count <= _T_27 ? _GEN_162 : L0Memory_33; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_263 = count >= 10'h1 & count <= _T_27 ? _GEN_163 : L0Memory_34; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_264 = count >= 10'h1 & count <= _T_27 ? _GEN_164 : L0Memory_35; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_265 = count >= 10'h1 & count <= _T_27 ? _GEN_165 : L0Memory_36; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_266 = count >= 10'h1 & count <= _T_27 ? _GEN_166 : L0Memory_37; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_267 = count >= 10'h1 & count <= _T_27 ? _GEN_167 : L0Memory_38; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_268 = count >= 10'h1 & count <= _T_27 ? _GEN_168 : L0Memory_39; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_269 = count >= 10'h1 & count <= _T_27 ? _GEN_169 : L0Memory_40; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_270 = count >= 10'h1 & count <= _T_27 ? _GEN_170 : L0Memory_41; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_271 = count >= 10'h1 & count <= _T_27 ? _GEN_171 : L0Memory_42; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_272 = count >= 10'h1 & count <= _T_27 ? _GEN_172 : L0Memory_43; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_273 = count >= 10'h1 & count <= _T_27 ? _GEN_173 : L0Memory_44; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_274 = count >= 10'h1 & count <= _T_27 ? _GEN_174 : L0Memory_45; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_275 = count >= 10'h1 & count <= _T_27 ? _GEN_175 : L0Memory_46; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_276 = count >= 10'h1 & count <= _T_27 ? _GEN_176 : L0Memory_47; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_277 = count >= 10'h1 & count <= _T_27 ? _GEN_177 : L0Memory_48; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_278 = count >= 10'h1 & count <= _T_27 ? _GEN_178 : L0Memory_49; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_279 = count >= 10'h1 & count <= _T_27 ? _GEN_179 : L0Memory_50; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_280 = count >= 10'h1 & count <= _T_27 ? _GEN_180 : L0Memory_51; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_281 = count >= 10'h1 & count <= _T_27 ? _GEN_181 : L0Memory_52; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_282 = count >= 10'h1 & count <= _T_27 ? _GEN_182 : L0Memory_53; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_283 = count >= 10'h1 & count <= _T_27 ? _GEN_183 : L0Memory_54; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_284 = count >= 10'h1 & count <= _T_27 ? _GEN_184 : L0Memory_55; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_285 = count >= 10'h1 & count <= _T_27 ? _GEN_185 : L0Memory_56; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_286 = count >= 10'h1 & count <= _T_27 ? _GEN_186 : L0Memory_57; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_287 = count >= 10'h1 & count <= _T_27 ? _GEN_187 : L0Memory_58; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_288 = count >= 10'h1 & count <= _T_27 ? _GEN_188 : L0Memory_59; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_289 = count >= 10'h1 & count <= _T_27 ? _GEN_189 : L0Memory_60; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_290 = count >= 10'h1 & count <= _T_27 ? _GEN_190 : L0Memory_61; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_291 = count >= 10'h1 & count <= _T_27 ? _GEN_191 : L0Memory_62; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_292 = count >= 10'h1 & count <= _T_27 ? _GEN_192 : L0Memory_63; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_293 = count >= 10'h1 & count <= _T_27 ? _GEN_193 : L0Memory_64; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_294 = count >= 10'h1 & count <= _T_27 ? _GEN_194 : L0Memory_65; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_295 = count >= 10'h1 & count <= _T_27 ? _GEN_195 : L0Memory_66; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_296 = count >= 10'h1 & count <= _T_27 ? _GEN_196 : L0Memory_67; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_297 = count >= 10'h1 & count <= _T_27 ? _GEN_197 : L0Memory_68; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_298 = count >= 10'h1 & count <= _T_27 ? _GEN_198 : L0Memory_69; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_299 = count >= 10'h1 & count <= _T_27 ? _GEN_199 : L0Memory_70; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_300 = count >= 10'h1 & count <= _T_27 ? _GEN_200 : L0Memory_71; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_301 = count >= 10'h1 & count <= _T_27 ? _GEN_201 : L0Memory_72; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_302 = count >= 10'h1 & count <= _T_27 ? _GEN_202 : L0Memory_73; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_303 = count >= 10'h1 & count <= _T_27 ? _GEN_203 : L0Memory_74; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_304 = count >= 10'h1 & count <= _T_27 ? _GEN_204 : L0Memory_75; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_305 = count >= 10'h1 & count <= _T_27 ? _GEN_205 : L0Memory_76; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_306 = count >= 10'h1 & count <= _T_27 ? _GEN_206 : L0Memory_77; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_307 = count >= 10'h1 & count <= _T_27 ? _GEN_207 : L0Memory_78; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_308 = count >= 10'h1 & count <= _T_27 ? _GEN_208 : L0Memory_79; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_309 = count >= 10'h1 & count <= _T_27 ? _GEN_209 : L0Memory_80; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_310 = count >= 10'h1 & count <= _T_27 ? _GEN_210 : L0Memory_81; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_311 = count >= 10'h1 & count <= _T_27 ? _GEN_211 : L0Memory_82; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_312 = count >= 10'h1 & count <= _T_27 ? _GEN_212 : L0Memory_83; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_313 = count >= 10'h1 & count <= _T_27 ? _GEN_213 : L0Memory_84; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_314 = count >= 10'h1 & count <= _T_27 ? _GEN_214 : L0Memory_85; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_315 = count >= 10'h1 & count <= _T_27 ? _GEN_215 : L0Memory_86; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_316 = count >= 10'h1 & count <= _T_27 ? _GEN_216 : L0Memory_87; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_317 = count >= 10'h1 & count <= _T_27 ? _GEN_217 : L0Memory_88; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_318 = count >= 10'h1 & count <= _T_27 ? _GEN_218 : L0Memory_89; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_319 = count >= 10'h1 & count <= _T_27 ? _GEN_219 : L0Memory_90; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_320 = count >= 10'h1 & count <= _T_27 ? _GEN_220 : L0Memory_91; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_321 = count >= 10'h1 & count <= _T_27 ? _GEN_221 : L0Memory_92; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_322 = count >= 10'h1 & count <= _T_27 ? _GEN_222 : L0Memory_93; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_323 = count >= 10'h1 & count <= _T_27 ? _GEN_223 : L0Memory_94; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_324 = count >= 10'h1 & count <= _T_27 ? _GEN_224 : L0Memory_95; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_325 = count >= 10'h1 & count <= _T_27 ? _GEN_225 : L0Memory_96; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_326 = count >= 10'h1 & count <= _T_27 ? _GEN_226 : L0Memory_97; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_327 = count >= 10'h1 & count <= _T_27 ? _GEN_227 : L0Memory_98; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_328 = count >= 10'h1 & count <= _T_27 ? _GEN_228 : L0Memory_99; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [5:0] _GEN_329 = count >= 10'h1 & count <= _T_27 ? _L0Index_T_2 : _GEN_128; // @[PEArray.scala 198:59 PEArray.scala 200:17]
  wire [9:0] _GEN_330 = _T_24 ? 10'h0 : _GEN_127; // @[PEArray.scala 202:32 PEArray.scala 203:15]
  wire [2:0] _GEN_331 = _T_24 ? 3'h0 : state; // @[PEArray.scala 202:32 PEArray.scala 204:15 PEArray.scala 100:22]
  wire [9:0] _GEN_865 = {{4'd0}, GRU_out_width}; // @[PEArray.scala 220:19]
  wire [9:0] _GEN_0 = count % _GEN_865; // @[PEArray.scala 220:19]
  wire [5:0] _T_36 = _GEN_0[5:0]; // @[PEArray.scala 220:19]
  wire [5:0] _T_38 = GRU_out_width - 6'h1; // @[PEArray.scala 220:55]
  wire [5:0] _GEN_334 = _T_36 == _T_38 ? _L0Index_T_2 : 6'h0; // @[PEArray.scala 220:62 PEArray.scala 221:17 PEArray.scala 214:15]
  wire [5:0] _GEN_346 = _T_41 ? _GEN_334 : L0Index; // @[Conditional.scala 39:67 PEArray.scala 39:24]
  wire [9:0] _GEN_347 = _T_41 ? _GEN_330 : count; // @[Conditional.scala 39:67 PEArray.scala 101:22]
  wire [2:0] _GEN_348 = _T_41 ? _GEN_331 : state; // @[Conditional.scala 39:67 PEArray.scala 100:22]
  wire [5:0] _GEN_353 = _T_31 ? _GEN_334 : _GEN_346; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_354 = _T_31 ? _GEN_330 : _GEN_347; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_355 = _T_31 ? _GEN_331 : _GEN_348; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_356 = _T_22 ? _GEN_330 : _GEN_354; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_357 = _T_22 ? _GEN_329 : _GEN_353; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_458 = _T_22 ? _GEN_331 : _GEN_355; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_690 = _T_3 ? _GEN_118 : {{2'd0}, GRU_out_width}; // @[Conditional.scala 40:58 PEArray.scala 104:26]
  FP16MulAdder FP16MAC ( // @[PEArray.scala 72:23]
    .io_a(FP16MAC_io_a),
    .io_b(FP16MAC_io_b),
    .io_c(FP16MAC_io_c),
    .io_out(FP16MAC_io_out)
  );
  assign io_ToRightPE = mux3out_reg; // @[PEArray.scala 95:16]
  assign io_ToBelowPE = mux2out_reg; // @[PEArray.scala 94:16]
  assign FP16MAC_io_a = sel1 ? io_FromL1 : io_FromLeftPE; // @[PEArray.scala 50:14 PEArray.scala 50:23 PEArray.scala 51:24]
  assign FP16MAC_io_b = sel5 ? mux4out : _GEN_105; // @[PEArray.scala 77:13 PEArray.scala 78:18 PEArray.scala 81:18]
  assign FP16MAC_io_c = sel5 ? _GEN_105 : mux4out; // @[PEArray.scala 77:13 PEArray.scala 79:18 PEArray.scala 82:18]
  always @(posedge clock) begin
    if (reset) begin // @[PEArray.scala 39:24]
      L0Index <= 6'h0; // @[PEArray.scala 39:24]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h1; // @[PEArray.scala 159:15]
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        L0Index <= 6'hb; // @[PEArray.scala 181:15]
      end else begin
        L0Index <= _GEN_357;
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_0 <= _GEN_229;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_1 <= _GEN_230;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_2 <= _GEN_231;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_3 <= _GEN_232;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_4 <= _GEN_233;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_5 <= _GEN_234;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_6 <= _GEN_235;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_7 <= _GEN_236;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_8 <= _GEN_237;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_9 <= _GEN_238;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_10 <= _GEN_239;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_11 <= _GEN_240;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_12 <= _GEN_241;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_13 <= _GEN_242;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_14 <= _GEN_243;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_15 <= _GEN_244;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_16 <= _GEN_245;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_17 <= _GEN_246;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_18 <= _GEN_247;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_19 <= _GEN_248;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_20 <= _GEN_249;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_21 <= _GEN_250;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_22 <= _GEN_251;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_23 <= _GEN_252;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_24 <= _GEN_253;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_25 <= _GEN_254;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_26 <= _GEN_255;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_27 <= _GEN_256;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_28 <= _GEN_257;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_29 <= _GEN_258;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_30 <= _GEN_259;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_31 <= _GEN_260;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_32 <= _GEN_261;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_33 <= _GEN_262;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_34 <= _GEN_263;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_35 <= _GEN_264;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_36 <= _GEN_265;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_37 <= _GEN_266;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_38 <= _GEN_267;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_39 <= _GEN_268;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_40 <= _GEN_269;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_41 <= _GEN_270;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_42 <= _GEN_271;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_43 <= _GEN_272;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_44 <= _GEN_273;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_45 <= _GEN_274;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_46 <= _GEN_275;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_47 <= _GEN_276;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_48 <= _GEN_277;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_49 <= _GEN_278;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_50 <= _GEN_279;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_51 <= _GEN_280;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_52 <= _GEN_281;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_53 <= _GEN_282;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_54 <= _GEN_283;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_55 <= _GEN_284;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_56 <= _GEN_285;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_57 <= _GEN_286;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_58 <= _GEN_287;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_59 <= _GEN_288;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_60 <= _GEN_289;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_61 <= _GEN_290;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_62 <= _GEN_291;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_63 <= _GEN_292;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_64 <= _GEN_293;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_65 <= _GEN_294;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_66 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_67 <= _GEN_296;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_68 <= _GEN_297;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_69 <= _GEN_298;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_70 <= _GEN_299;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_71 <= _GEN_300;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_72 <= _GEN_301;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_73 <= _GEN_302;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_74 <= _GEN_303;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_75 <= _GEN_304;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_76 <= _GEN_305;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_77 <= _GEN_306;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_78 <= _GEN_307;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_79 <= _GEN_308;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_80 <= _GEN_309;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_81 <= _GEN_310;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_82 <= _GEN_311;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_83 <= _GEN_312;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_84 <= _GEN_313;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_85 <= _GEN_314;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_86 <= _GEN_315;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_87 <= _GEN_316;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_88 <= _GEN_317;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_89 <= _GEN_318;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_90 <= _GEN_319;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_91 <= _GEN_320;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_92 <= _GEN_321;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_93 <= _GEN_322;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_94 <= _GEN_323;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_95 <= _GEN_324;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_96 <= _GEN_325;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_97 <= _GEN_326;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_98 <= _GEN_327;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_99 <= _GEN_328;
          end
        end
      end
    end
    if (reset) begin // @[PEArray.scala 100:22]
      state <= 3'h0; // @[PEArray.scala 100:22]
    end else if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[3]) begin // @[PEArray.scala 116:57]
        state <= 3'h1;
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      if (count == 10'h33) begin // @[PEArray.scala 164:27]
        state <= 3'h0; // @[PEArray.scala 166:15]
      end
    end else if (_T_16) begin // @[Conditional.scala 39:67]
      state <= _GEN_126;
    end else begin
      state <= _GEN_458;
    end
    if (reset) begin // @[PEArray.scala 90:28]
      mux2out_reg <= 16'h0; // @[PEArray.scala 90:28]
    end else begin
      mux2out_reg <= MAC_out; // @[PEArray.scala 90:28]
    end
    if (reset) begin // @[PEArray.scala 91:28]
      mux3out_reg <= 16'h0; // @[PEArray.scala 91:28]
    end else if (sel3) begin // @[PEArray.scala 56:14]
      mux3out_reg <= MAC_out; // @[PEArray.scala 56:23]
    end else if (sel1) begin // @[PEArray.scala 50:14]
      mux3out_reg <= io_FromL1; // @[PEArray.scala 50:23]
    end else begin
      mux3out_reg <= io_FromLeftPE; // @[PEArray.scala 51:24]
    end
    if (reset) begin // @[PEArray.scala 101:22]
      count <= 10'h0; // @[PEArray.scala 101:22]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        if (count == 10'h33) begin // @[PEArray.scala 164:27]
          count <= 10'h0; // @[PEArray.scala 165:15]
        end else begin
          count <= _GEN_120;
        end
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        count <= _GEN_125;
      end else begin
        count <= _GEN_356;
      end
    end
    GRU_out_width <= _GEN_690[5:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  L0Index = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  L0Memory_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  L0Memory_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  L0Memory_2 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  L0Memory_3 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  L0Memory_4 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  L0Memory_5 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  L0Memory_6 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  L0Memory_7 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  L0Memory_8 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  L0Memory_9 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  L0Memory_10 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  L0Memory_11 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  L0Memory_12 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  L0Memory_13 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  L0Memory_14 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  L0Memory_15 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  L0Memory_16 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  L0Memory_17 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  L0Memory_18 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  L0Memory_19 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  L0Memory_20 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  L0Memory_21 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  L0Memory_22 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  L0Memory_23 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  L0Memory_24 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  L0Memory_25 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  L0Memory_26 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  L0Memory_27 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  L0Memory_28 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  L0Memory_29 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  L0Memory_30 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  L0Memory_31 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  L0Memory_32 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  L0Memory_33 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  L0Memory_34 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  L0Memory_35 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  L0Memory_36 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  L0Memory_37 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  L0Memory_38 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  L0Memory_39 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  L0Memory_40 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  L0Memory_41 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  L0Memory_42 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  L0Memory_43 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  L0Memory_44 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  L0Memory_45 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  L0Memory_46 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  L0Memory_47 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  L0Memory_48 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  L0Memory_49 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  L0Memory_50 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  L0Memory_51 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  L0Memory_52 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  L0Memory_53 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  L0Memory_54 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  L0Memory_55 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  L0Memory_56 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  L0Memory_57 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  L0Memory_58 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  L0Memory_59 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  L0Memory_60 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  L0Memory_61 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  L0Memory_62 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  L0Memory_63 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  L0Memory_64 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  L0Memory_65 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  L0Memory_66 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  L0Memory_67 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  L0Memory_68 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  L0Memory_69 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  L0Memory_70 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  L0Memory_71 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  L0Memory_72 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  L0Memory_73 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  L0Memory_74 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  L0Memory_75 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  L0Memory_76 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  L0Memory_77 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  L0Memory_78 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  L0Memory_79 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  L0Memory_80 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  L0Memory_81 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  L0Memory_82 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  L0Memory_83 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  L0Memory_84 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  L0Memory_85 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  L0Memory_86 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  L0Memory_87 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  L0Memory_88 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  L0Memory_89 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  L0Memory_90 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  L0Memory_91 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  L0Memory_92 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  L0Memory_93 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  L0Memory_94 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  L0Memory_95 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  L0Memory_96 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  L0Memory_97 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  L0Memory_98 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  L0Memory_99 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  state = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  mux2out_reg = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  mux3out_reg = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  count = _RAND_104[9:0];
  _RAND_105 = {1{`RANDOM}};
  GRU_out_width = _RAND_105[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PE_26(
  input         clock,
  input         reset,
  input  [15:0] io_FromAbovePE,
  input  [15:0] io_FromLeftPE,
  input  [15:0] io_FromL1,
  input  [2:0]  io_control_signal_control,
  input  [9:0]  io_control_signal_count,
  input  [5:0]  io_control_signal_L0index,
  input  [11:0] io_control_signal_mask,
  input  [7:0]  io_control_signal_gru_out_width,
  output [15:0] io_ToRightPE,
  output [15:0] io_ToBelowPE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] FP16MAC_io_a; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_b; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_c; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_out; // @[PEArray.scala 72:23]
  reg [5:0] L0Index; // @[PEArray.scala 39:24]
  reg [15:0] L0Memory_0; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_1; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_2; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_3; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_4; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_5; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_6; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_7; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_8; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_9; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_10; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_11; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_12; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_13; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_14; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_15; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_16; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_17; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_18; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_19; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_20; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_21; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_22; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_23; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_24; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_25; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_26; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_27; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_28; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_29; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_30; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_31; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_32; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_33; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_34; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_35; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_36; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_37; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_38; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_39; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_40; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_41; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_42; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_43; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_44; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_45; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_46; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_47; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_48; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_49; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_50; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_51; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_52; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_53; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_54; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_55; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_56; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_57; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_58; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_59; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_60; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_61; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_62; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_63; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_64; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_65; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_66; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_67; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_68; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_69; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_70; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_71; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_72; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_73; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_74; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_75; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_76; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_77; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_78; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_79; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_80; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_81; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_82; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_83; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_84; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_85; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_86; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_87; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_88; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_89; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_90; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_91; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_92; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_93; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_94; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_95; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_96; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_97; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_98; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_99; // @[PEArray.scala 40:21]
  reg [2:0] state; // @[PEArray.scala 100:22]
  wire  _T_3 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_12 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_16 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_22 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_31 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_41 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_342 = _T_41 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 231:12 PEArray.scala 32:8]
  wire  _GEN_349 = _T_31 ? 1'h0 : _GEN_342; // @[Conditional.scala 39:67 PEArray.scala 208:12]
  wire  _GEN_459 = _T_22 | _GEN_349; // @[Conditional.scala 39:67 PEArray.scala 32:8]
  wire  _GEN_463 = _T_16 ? 1'h0 : _GEN_459; // @[Conditional.scala 39:67]
  wire  _GEN_572 = _T_12 | _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 149:12]
  wire  sel1 = _T_3 | _GEN_572; // @[Conditional.scala 40:58 PEArray.scala 108:12]
  wire [15:0] MAC_out = FP16MAC_io_out; // @[PEArray.scala 47:21 PEArray.scala 85:11]
  wire  _GEN_465 = _T_16 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 177:12]
  wire  _GEN_580 = _T_12 | _GEN_465; // @[Conditional.scala 39:67 PEArray.scala 34:8]
  wire  sel3 = _T_3 | _GEN_580; // @[Conditional.scala 40:58 PEArray.scala 110:12]
  wire [1:0] _GEN_344 = _T_41 ? 2'h2 : 2'h0; // @[Conditional.scala 39:67 PEArray.scala 233:12 PEArray.scala 35:8]
  wire [1:0] _GEN_351 = _T_31 ? 2'h2 : _GEN_344; // @[Conditional.scala 39:67 PEArray.scala 210:12]
  wire [1:0] _GEN_461 = _T_22 ? 2'h0 : _GEN_351; // @[Conditional.scala 39:67 PEArray.scala 35:8]
  wire [1:0] _GEN_466 = _T_16 ? 2'h0 : _GEN_461; // @[Conditional.scala 39:67 PEArray.scala 178:12]
  wire [1:0] _GEN_574 = _T_12 ? 2'h1 : _GEN_466; // @[Conditional.scala 39:67]
  wire [1:0] sel4 = _T_3 ? 2'h0 : _GEN_574; // @[Conditional.scala 40:58 PEArray.scala 111:12]
  wire [15:0] _GEN_3 = sel4 == 2'h2 ? io_FromL1 : 16'h0; // @[PEArray.scala 65:28 PEArray.scala 66:15 PEArray.scala 69:15]
  wire [15:0] _GEN_4 = sel4 == 2'h1 ? io_FromAbovePE : _GEN_3; // @[PEArray.scala 62:28 PEArray.scala 63:15]
  wire [15:0] mux4out = sel4 == 2'h0 ? 16'h0 : _GEN_4; // @[PEArray.scala 59:22 PEArray.scala 60:13]
  wire [15:0] _GEN_7 = 6'h1 == L0Index ? L0Memory_1 : L0Memory_0; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_8 = 6'h2 == L0Index ? L0Memory_2 : _GEN_7; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_9 = 6'h3 == L0Index ? L0Memory_3 : _GEN_8; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_10 = 6'h4 == L0Index ? L0Memory_4 : _GEN_9; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_11 = 6'h5 == L0Index ? L0Memory_5 : _GEN_10; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_12 = 6'h6 == L0Index ? L0Memory_6 : _GEN_11; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_13 = 6'h7 == L0Index ? L0Memory_7 : _GEN_12; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_14 = 6'h8 == L0Index ? L0Memory_8 : _GEN_13; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_15 = 6'h9 == L0Index ? L0Memory_9 : _GEN_14; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_16 = 6'ha == L0Index ? L0Memory_10 : _GEN_15; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_17 = 6'hb == L0Index ? L0Memory_11 : _GEN_16; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_18 = 6'hc == L0Index ? L0Memory_12 : _GEN_17; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_19 = 6'hd == L0Index ? L0Memory_13 : _GEN_18; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_20 = 6'he == L0Index ? L0Memory_14 : _GEN_19; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_21 = 6'hf == L0Index ? L0Memory_15 : _GEN_20; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_22 = 6'h10 == L0Index ? L0Memory_16 : _GEN_21; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_23 = 6'h11 == L0Index ? L0Memory_17 : _GEN_22; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_24 = 6'h12 == L0Index ? L0Memory_18 : _GEN_23; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_25 = 6'h13 == L0Index ? L0Memory_19 : _GEN_24; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_26 = 6'h14 == L0Index ? L0Memory_20 : _GEN_25; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_27 = 6'h15 == L0Index ? L0Memory_21 : _GEN_26; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_28 = 6'h16 == L0Index ? L0Memory_22 : _GEN_27; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_29 = 6'h17 == L0Index ? L0Memory_23 : _GEN_28; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_30 = 6'h18 == L0Index ? L0Memory_24 : _GEN_29; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_31 = 6'h19 == L0Index ? L0Memory_25 : _GEN_30; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_32 = 6'h1a == L0Index ? L0Memory_26 : _GEN_31; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_33 = 6'h1b == L0Index ? L0Memory_27 : _GEN_32; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_34 = 6'h1c == L0Index ? L0Memory_28 : _GEN_33; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_35 = 6'h1d == L0Index ? L0Memory_29 : _GEN_34; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_36 = 6'h1e == L0Index ? L0Memory_30 : _GEN_35; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_37 = 6'h1f == L0Index ? L0Memory_31 : _GEN_36; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_38 = 6'h20 == L0Index ? L0Memory_32 : _GEN_37; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_39 = 6'h21 == L0Index ? L0Memory_33 : _GEN_38; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_40 = 6'h22 == L0Index ? L0Memory_34 : _GEN_39; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_41 = 6'h23 == L0Index ? L0Memory_35 : _GEN_40; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_42 = 6'h24 == L0Index ? L0Memory_36 : _GEN_41; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_43 = 6'h25 == L0Index ? L0Memory_37 : _GEN_42; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_44 = 6'h26 == L0Index ? L0Memory_38 : _GEN_43; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_45 = 6'h27 == L0Index ? L0Memory_39 : _GEN_44; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_46 = 6'h28 == L0Index ? L0Memory_40 : _GEN_45; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_47 = 6'h29 == L0Index ? L0Memory_41 : _GEN_46; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_48 = 6'h2a == L0Index ? L0Memory_42 : _GEN_47; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_49 = 6'h2b == L0Index ? L0Memory_43 : _GEN_48; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_50 = 6'h2c == L0Index ? L0Memory_44 : _GEN_49; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_51 = 6'h2d == L0Index ? L0Memory_45 : _GEN_50; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_52 = 6'h2e == L0Index ? L0Memory_46 : _GEN_51; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_53 = 6'h2f == L0Index ? L0Memory_47 : _GEN_52; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_54 = 6'h30 == L0Index ? L0Memory_48 : _GEN_53; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_55 = 6'h31 == L0Index ? L0Memory_49 : _GEN_54; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_56 = 6'h32 == L0Index ? L0Memory_50 : _GEN_55; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_57 = 6'h33 == L0Index ? L0Memory_51 : _GEN_56; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_58 = 6'h34 == L0Index ? L0Memory_52 : _GEN_57; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_59 = 6'h35 == L0Index ? L0Memory_53 : _GEN_58; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_60 = 6'h36 == L0Index ? L0Memory_54 : _GEN_59; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_61 = 6'h37 == L0Index ? L0Memory_55 : _GEN_60; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_62 = 6'h38 == L0Index ? L0Memory_56 : _GEN_61; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_63 = 6'h39 == L0Index ? L0Memory_57 : _GEN_62; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_64 = 6'h3a == L0Index ? L0Memory_58 : _GEN_63; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_65 = 6'h3b == L0Index ? L0Memory_59 : _GEN_64; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_66 = 6'h3c == L0Index ? L0Memory_60 : _GEN_65; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_67 = 6'h3d == L0Index ? L0Memory_61 : _GEN_66; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_68 = 6'h3e == L0Index ? L0Memory_62 : _GEN_67; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_69 = 6'h3f == L0Index ? L0Memory_63 : _GEN_68; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [6:0] _GEN_793 = {{1'd0}, L0Index}; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_70 = 7'h40 == _GEN_793 ? L0Memory_64 : _GEN_69; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_71 = 7'h41 == _GEN_793 ? L0Memory_65 : _GEN_70; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_72 = 7'h42 == _GEN_793 ? L0Memory_66 : _GEN_71; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_73 = 7'h43 == _GEN_793 ? L0Memory_67 : _GEN_72; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_74 = 7'h44 == _GEN_793 ? L0Memory_68 : _GEN_73; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_75 = 7'h45 == _GEN_793 ? L0Memory_69 : _GEN_74; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_76 = 7'h46 == _GEN_793 ? L0Memory_70 : _GEN_75; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_77 = 7'h47 == _GEN_793 ? L0Memory_71 : _GEN_76; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_78 = 7'h48 == _GEN_793 ? L0Memory_72 : _GEN_77; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_79 = 7'h49 == _GEN_793 ? L0Memory_73 : _GEN_78; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_80 = 7'h4a == _GEN_793 ? L0Memory_74 : _GEN_79; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_81 = 7'h4b == _GEN_793 ? L0Memory_75 : _GEN_80; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_82 = 7'h4c == _GEN_793 ? L0Memory_76 : _GEN_81; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_83 = 7'h4d == _GEN_793 ? L0Memory_77 : _GEN_82; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_84 = 7'h4e == _GEN_793 ? L0Memory_78 : _GEN_83; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_85 = 7'h4f == _GEN_793 ? L0Memory_79 : _GEN_84; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_86 = 7'h50 == _GEN_793 ? L0Memory_80 : _GEN_85; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_87 = 7'h51 == _GEN_793 ? L0Memory_81 : _GEN_86; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_88 = 7'h52 == _GEN_793 ? L0Memory_82 : _GEN_87; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_89 = 7'h53 == _GEN_793 ? L0Memory_83 : _GEN_88; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_90 = 7'h54 == _GEN_793 ? L0Memory_84 : _GEN_89; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_91 = 7'h55 == _GEN_793 ? L0Memory_85 : _GEN_90; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_92 = 7'h56 == _GEN_793 ? L0Memory_86 : _GEN_91; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_93 = 7'h57 == _GEN_793 ? L0Memory_87 : _GEN_92; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_94 = 7'h58 == _GEN_793 ? L0Memory_88 : _GEN_93; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_95 = 7'h59 == _GEN_793 ? L0Memory_89 : _GEN_94; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_96 = 7'h5a == _GEN_793 ? L0Memory_90 : _GEN_95; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_97 = 7'h5b == _GEN_793 ? L0Memory_91 : _GEN_96; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_98 = 7'h5c == _GEN_793 ? L0Memory_92 : _GEN_97; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_99 = 7'h5d == _GEN_793 ? L0Memory_93 : _GEN_98; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_100 = 7'h5e == _GEN_793 ? L0Memory_94 : _GEN_99; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_101 = 7'h5f == _GEN_793 ? L0Memory_95 : _GEN_100; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_102 = 7'h60 == _GEN_793 ? L0Memory_96 : _GEN_101; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_103 = 7'h61 == _GEN_793 ? L0Memory_97 : _GEN_102; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_104 = 7'h62 == _GEN_793 ? L0Memory_98 : _GEN_103; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_105 = 7'h63 == _GEN_793 ? L0Memory_99 : _GEN_104; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire  _GEN_575 = _T_12 ? 1'h0 : _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 157:12]
  wire  sel5 = _T_3 ? 1'h0 : _GEN_575; // @[Conditional.scala 40:58 PEArray.scala 112:12]
  reg [15:0] mux2out_reg; // @[PEArray.scala 90:28]
  reg [15:0] mux3out_reg; // @[PEArray.scala 91:28]
  reg [9:0] count; // @[PEArray.scala 101:22]
  reg [9:0] count_max; // @[PEArray.scala 102:22]
  reg [5:0] L0index_begin; // @[PEArray.scala 103:26]
  reg [5:0] GRU_out_width; // @[PEArray.scala 104:26]
  wire  _T_6 = 3'h0 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_7 = 3'h1 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_8 = 3'h2 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_9 = 3'h3 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_10 = 3'h4 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_11 = 3'h5 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_109 = _T_11 ? 3'h5 : state; // @[Conditional.scala 39:67 PEArray.scala 140:19 PEArray.scala 100:22]
  wire [2:0] _GEN_110 = _T_10 ? 3'h4 : _GEN_109; // @[Conditional.scala 39:67 PEArray.scala 136:19]
  wire [2:0] _GEN_111 = _T_9 ? 3'h3 : _GEN_110; // @[Conditional.scala 39:67 PEArray.scala 132:19]
  wire [2:0] _GEN_112 = _T_8 ? 3'h2 : _GEN_111; // @[Conditional.scala 39:67 PEArray.scala 128:19]
  wire [2:0] _GEN_113 = _T_7 ? 3'h1 : _GEN_112; // @[Conditional.scala 39:67 PEArray.scala 124:19]
  wire [7:0] _GEN_118 = io_control_signal_mask[3] ? io_control_signal_gru_out_width : {{2'd0}, GRU_out_width}; // @[PEArray.scala 116:57 PEArray.scala 145:23 PEArray.scala 104:26]
  wire [9:0] _count_T_1 = count + 10'h1; // @[PEArray.scala 162:24]
  wire [9:0] _GEN_120 = count != 10'h33 ? _count_T_1 : count; // @[PEArray.scala 161:27 PEArray.scala 162:15 PEArray.scala 101:22]
  wire [9:0] _GEN_124 = count != 10'h188 ? _count_T_1 : count; // @[PEArray.scala 183:28 PEArray.scala 184:15 PEArray.scala 101:22]
  wire [9:0] _GEN_125 = count == 10'h188 ? 10'h0 : _GEN_124; // @[PEArray.scala 186:28 PEArray.scala 187:15]
  wire [2:0] _GEN_126 = count == 10'h188 ? 3'h0 : state; // @[PEArray.scala 186:28 PEArray.scala 188:15 PEArray.scala 100:22]
  wire [9:0] _GEN_127 = count != count_max ? _count_T_1 : count; // @[PEArray.scala 192:32 PEArray.scala 193:15 PEArray.scala 101:22]
  wire [5:0] _GEN_128 = count == 10'h0 ? L0index_begin : L0Index; // @[PEArray.scala 195:26 PEArray.scala 196:17 PEArray.scala 39:24]
  wire [9:0] _T_27 = count_max - 10'h1; // @[PEArray.scala 198:51]
  wire [15:0] _GEN_129 = 6'h0 == L0Index ? io_FromL1 : L0Memory_0; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_130 = 6'h1 == L0Index ? io_FromL1 : L0Memory_1; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_131 = 6'h2 == L0Index ? io_FromL1 : L0Memory_2; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_132 = 6'h3 == L0Index ? io_FromL1 : L0Memory_3; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_133 = 6'h4 == L0Index ? io_FromL1 : L0Memory_4; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_134 = 6'h5 == L0Index ? io_FromL1 : L0Memory_5; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_135 = 6'h6 == L0Index ? io_FromL1 : L0Memory_6; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_136 = 6'h7 == L0Index ? io_FromL1 : L0Memory_7; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_137 = 6'h8 == L0Index ? io_FromL1 : L0Memory_8; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_138 = 6'h9 == L0Index ? io_FromL1 : L0Memory_9; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_139 = 6'ha == L0Index ? io_FromL1 : L0Memory_10; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_140 = 6'hb == L0Index ? io_FromL1 : L0Memory_11; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_141 = 6'hc == L0Index ? io_FromL1 : L0Memory_12; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_142 = 6'hd == L0Index ? io_FromL1 : L0Memory_13; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_143 = 6'he == L0Index ? io_FromL1 : L0Memory_14; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_144 = 6'hf == L0Index ? io_FromL1 : L0Memory_15; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_145 = 6'h10 == L0Index ? io_FromL1 : L0Memory_16; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_146 = 6'h11 == L0Index ? io_FromL1 : L0Memory_17; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_147 = 6'h12 == L0Index ? io_FromL1 : L0Memory_18; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_148 = 6'h13 == L0Index ? io_FromL1 : L0Memory_19; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_149 = 6'h14 == L0Index ? io_FromL1 : L0Memory_20; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_150 = 6'h15 == L0Index ? io_FromL1 : L0Memory_21; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_151 = 6'h16 == L0Index ? io_FromL1 : L0Memory_22; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_152 = 6'h17 == L0Index ? io_FromL1 : L0Memory_23; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_153 = 6'h18 == L0Index ? io_FromL1 : L0Memory_24; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_154 = 6'h19 == L0Index ? io_FromL1 : L0Memory_25; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_155 = 6'h1a == L0Index ? io_FromL1 : L0Memory_26; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_156 = 6'h1b == L0Index ? io_FromL1 : L0Memory_27; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_157 = 6'h1c == L0Index ? io_FromL1 : L0Memory_28; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_158 = 6'h1d == L0Index ? io_FromL1 : L0Memory_29; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_159 = 6'h1e == L0Index ? io_FromL1 : L0Memory_30; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_160 = 6'h1f == L0Index ? io_FromL1 : L0Memory_31; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_161 = 6'h20 == L0Index ? io_FromL1 : L0Memory_32; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_162 = 6'h21 == L0Index ? io_FromL1 : L0Memory_33; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_163 = 6'h22 == L0Index ? io_FromL1 : L0Memory_34; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_164 = 6'h23 == L0Index ? io_FromL1 : L0Memory_35; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_165 = 6'h24 == L0Index ? io_FromL1 : L0Memory_36; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_166 = 6'h25 == L0Index ? io_FromL1 : L0Memory_37; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_167 = 6'h26 == L0Index ? io_FromL1 : L0Memory_38; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_168 = 6'h27 == L0Index ? io_FromL1 : L0Memory_39; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_169 = 6'h28 == L0Index ? io_FromL1 : L0Memory_40; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_170 = 6'h29 == L0Index ? io_FromL1 : L0Memory_41; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_171 = 6'h2a == L0Index ? io_FromL1 : L0Memory_42; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_172 = 6'h2b == L0Index ? io_FromL1 : L0Memory_43; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_173 = 6'h2c == L0Index ? io_FromL1 : L0Memory_44; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_174 = 6'h2d == L0Index ? io_FromL1 : L0Memory_45; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_175 = 6'h2e == L0Index ? io_FromL1 : L0Memory_46; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_176 = 6'h2f == L0Index ? io_FromL1 : L0Memory_47; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_177 = 6'h30 == L0Index ? io_FromL1 : L0Memory_48; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_178 = 6'h31 == L0Index ? io_FromL1 : L0Memory_49; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_179 = 6'h32 == L0Index ? io_FromL1 : L0Memory_50; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_180 = 6'h33 == L0Index ? io_FromL1 : L0Memory_51; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_181 = 6'h34 == L0Index ? io_FromL1 : L0Memory_52; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_182 = 6'h35 == L0Index ? io_FromL1 : L0Memory_53; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_183 = 6'h36 == L0Index ? io_FromL1 : L0Memory_54; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_184 = 6'h37 == L0Index ? io_FromL1 : L0Memory_55; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_185 = 6'h38 == L0Index ? io_FromL1 : L0Memory_56; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_186 = 6'h39 == L0Index ? io_FromL1 : L0Memory_57; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_187 = 6'h3a == L0Index ? io_FromL1 : L0Memory_58; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_188 = 6'h3b == L0Index ? io_FromL1 : L0Memory_59; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_189 = 6'h3c == L0Index ? io_FromL1 : L0Memory_60; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_190 = 6'h3d == L0Index ? io_FromL1 : L0Memory_61; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_191 = 6'h3e == L0Index ? io_FromL1 : L0Memory_62; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_192 = 6'h3f == L0Index ? io_FromL1 : L0Memory_63; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_193 = 7'h40 == _GEN_793 ? io_FromL1 : L0Memory_64; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_194 = 7'h41 == _GEN_793 ? io_FromL1 : L0Memory_65; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_195 = 7'h42 == _GEN_793 ? io_FromL1 : L0Memory_66; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_196 = 7'h43 == _GEN_793 ? io_FromL1 : L0Memory_67; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_197 = 7'h44 == _GEN_793 ? io_FromL1 : L0Memory_68; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_198 = 7'h45 == _GEN_793 ? io_FromL1 : L0Memory_69; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_199 = 7'h46 == _GEN_793 ? io_FromL1 : L0Memory_70; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_200 = 7'h47 == _GEN_793 ? io_FromL1 : L0Memory_71; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_201 = 7'h48 == _GEN_793 ? io_FromL1 : L0Memory_72; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_202 = 7'h49 == _GEN_793 ? io_FromL1 : L0Memory_73; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_203 = 7'h4a == _GEN_793 ? io_FromL1 : L0Memory_74; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_204 = 7'h4b == _GEN_793 ? io_FromL1 : L0Memory_75; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_205 = 7'h4c == _GEN_793 ? io_FromL1 : L0Memory_76; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_206 = 7'h4d == _GEN_793 ? io_FromL1 : L0Memory_77; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_207 = 7'h4e == _GEN_793 ? io_FromL1 : L0Memory_78; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_208 = 7'h4f == _GEN_793 ? io_FromL1 : L0Memory_79; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_209 = 7'h50 == _GEN_793 ? io_FromL1 : L0Memory_80; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_210 = 7'h51 == _GEN_793 ? io_FromL1 : L0Memory_81; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_211 = 7'h52 == _GEN_793 ? io_FromL1 : L0Memory_82; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_212 = 7'h53 == _GEN_793 ? io_FromL1 : L0Memory_83; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_213 = 7'h54 == _GEN_793 ? io_FromL1 : L0Memory_84; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_214 = 7'h55 == _GEN_793 ? io_FromL1 : L0Memory_85; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_215 = 7'h56 == _GEN_793 ? io_FromL1 : L0Memory_86; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_216 = 7'h57 == _GEN_793 ? io_FromL1 : L0Memory_87; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_217 = 7'h58 == _GEN_793 ? io_FromL1 : L0Memory_88; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_218 = 7'h59 == _GEN_793 ? io_FromL1 : L0Memory_89; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_219 = 7'h5a == _GEN_793 ? io_FromL1 : L0Memory_90; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_220 = 7'h5b == _GEN_793 ? io_FromL1 : L0Memory_91; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_221 = 7'h5c == _GEN_793 ? io_FromL1 : L0Memory_92; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_222 = 7'h5d == _GEN_793 ? io_FromL1 : L0Memory_93; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_223 = 7'h5e == _GEN_793 ? io_FromL1 : L0Memory_94; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_224 = 7'h5f == _GEN_793 ? io_FromL1 : L0Memory_95; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_225 = 7'h60 == _GEN_793 ? io_FromL1 : L0Memory_96; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_226 = 7'h61 == _GEN_793 ? io_FromL1 : L0Memory_97; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_227 = 7'h62 == _GEN_793 ? io_FromL1 : L0Memory_98; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_228 = 7'h63 == _GEN_793 ? io_FromL1 : L0Memory_99; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [5:0] _L0Index_T_2 = L0Index + 6'h1; // @[PEArray.scala 200:28]
  wire [15:0] _GEN_229 = count >= 10'h1 & count <= _T_27 ? _GEN_129 : L0Memory_0; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_230 = count >= 10'h1 & count <= _T_27 ? _GEN_130 : L0Memory_1; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_231 = count >= 10'h1 & count <= _T_27 ? _GEN_131 : L0Memory_2; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_232 = count >= 10'h1 & count <= _T_27 ? _GEN_132 : L0Memory_3; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_233 = count >= 10'h1 & count <= _T_27 ? _GEN_133 : L0Memory_4; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_234 = count >= 10'h1 & count <= _T_27 ? _GEN_134 : L0Memory_5; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_235 = count >= 10'h1 & count <= _T_27 ? _GEN_135 : L0Memory_6; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_236 = count >= 10'h1 & count <= _T_27 ? _GEN_136 : L0Memory_7; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_237 = count >= 10'h1 & count <= _T_27 ? _GEN_137 : L0Memory_8; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_238 = count >= 10'h1 & count <= _T_27 ? _GEN_138 : L0Memory_9; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_239 = count >= 10'h1 & count <= _T_27 ? _GEN_139 : L0Memory_10; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_240 = count >= 10'h1 & count <= _T_27 ? _GEN_140 : L0Memory_11; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_241 = count >= 10'h1 & count <= _T_27 ? _GEN_141 : L0Memory_12; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_242 = count >= 10'h1 & count <= _T_27 ? _GEN_142 : L0Memory_13; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_243 = count >= 10'h1 & count <= _T_27 ? _GEN_143 : L0Memory_14; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_244 = count >= 10'h1 & count <= _T_27 ? _GEN_144 : L0Memory_15; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_245 = count >= 10'h1 & count <= _T_27 ? _GEN_145 : L0Memory_16; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_246 = count >= 10'h1 & count <= _T_27 ? _GEN_146 : L0Memory_17; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_247 = count >= 10'h1 & count <= _T_27 ? _GEN_147 : L0Memory_18; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_248 = count >= 10'h1 & count <= _T_27 ? _GEN_148 : L0Memory_19; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_249 = count >= 10'h1 & count <= _T_27 ? _GEN_149 : L0Memory_20; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_250 = count >= 10'h1 & count <= _T_27 ? _GEN_150 : L0Memory_21; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_251 = count >= 10'h1 & count <= _T_27 ? _GEN_151 : L0Memory_22; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_252 = count >= 10'h1 & count <= _T_27 ? _GEN_152 : L0Memory_23; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_253 = count >= 10'h1 & count <= _T_27 ? _GEN_153 : L0Memory_24; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_254 = count >= 10'h1 & count <= _T_27 ? _GEN_154 : L0Memory_25; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_255 = count >= 10'h1 & count <= _T_27 ? _GEN_155 : L0Memory_26; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_256 = count >= 10'h1 & count <= _T_27 ? _GEN_156 : L0Memory_27; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_257 = count >= 10'h1 & count <= _T_27 ? _GEN_157 : L0Memory_28; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_258 = count >= 10'h1 & count <= _T_27 ? _GEN_158 : L0Memory_29; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_259 = count >= 10'h1 & count <= _T_27 ? _GEN_159 : L0Memory_30; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_260 = count >= 10'h1 & count <= _T_27 ? _GEN_160 : L0Memory_31; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_261 = count >= 10'h1 & count <= _T_27 ? _GEN_161 : L0Memory_32; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_262 = count >= 10'h1 & count <= _T_27 ? _GEN_162 : L0Memory_33; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_263 = count >= 10'h1 & count <= _T_27 ? _GEN_163 : L0Memory_34; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_264 = count >= 10'h1 & count <= _T_27 ? _GEN_164 : L0Memory_35; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_265 = count >= 10'h1 & count <= _T_27 ? _GEN_165 : L0Memory_36; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_266 = count >= 10'h1 & count <= _T_27 ? _GEN_166 : L0Memory_37; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_267 = count >= 10'h1 & count <= _T_27 ? _GEN_167 : L0Memory_38; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_268 = count >= 10'h1 & count <= _T_27 ? _GEN_168 : L0Memory_39; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_269 = count >= 10'h1 & count <= _T_27 ? _GEN_169 : L0Memory_40; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_270 = count >= 10'h1 & count <= _T_27 ? _GEN_170 : L0Memory_41; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_271 = count >= 10'h1 & count <= _T_27 ? _GEN_171 : L0Memory_42; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_272 = count >= 10'h1 & count <= _T_27 ? _GEN_172 : L0Memory_43; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_273 = count >= 10'h1 & count <= _T_27 ? _GEN_173 : L0Memory_44; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_274 = count >= 10'h1 & count <= _T_27 ? _GEN_174 : L0Memory_45; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_275 = count >= 10'h1 & count <= _T_27 ? _GEN_175 : L0Memory_46; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_276 = count >= 10'h1 & count <= _T_27 ? _GEN_176 : L0Memory_47; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_277 = count >= 10'h1 & count <= _T_27 ? _GEN_177 : L0Memory_48; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_278 = count >= 10'h1 & count <= _T_27 ? _GEN_178 : L0Memory_49; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_279 = count >= 10'h1 & count <= _T_27 ? _GEN_179 : L0Memory_50; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_280 = count >= 10'h1 & count <= _T_27 ? _GEN_180 : L0Memory_51; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_281 = count >= 10'h1 & count <= _T_27 ? _GEN_181 : L0Memory_52; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_282 = count >= 10'h1 & count <= _T_27 ? _GEN_182 : L0Memory_53; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_283 = count >= 10'h1 & count <= _T_27 ? _GEN_183 : L0Memory_54; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_284 = count >= 10'h1 & count <= _T_27 ? _GEN_184 : L0Memory_55; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_285 = count >= 10'h1 & count <= _T_27 ? _GEN_185 : L0Memory_56; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_286 = count >= 10'h1 & count <= _T_27 ? _GEN_186 : L0Memory_57; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_287 = count >= 10'h1 & count <= _T_27 ? _GEN_187 : L0Memory_58; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_288 = count >= 10'h1 & count <= _T_27 ? _GEN_188 : L0Memory_59; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_289 = count >= 10'h1 & count <= _T_27 ? _GEN_189 : L0Memory_60; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_290 = count >= 10'h1 & count <= _T_27 ? _GEN_190 : L0Memory_61; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_291 = count >= 10'h1 & count <= _T_27 ? _GEN_191 : L0Memory_62; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_292 = count >= 10'h1 & count <= _T_27 ? _GEN_192 : L0Memory_63; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_293 = count >= 10'h1 & count <= _T_27 ? _GEN_193 : L0Memory_64; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_294 = count >= 10'h1 & count <= _T_27 ? _GEN_194 : L0Memory_65; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_295 = count >= 10'h1 & count <= _T_27 ? _GEN_195 : L0Memory_66; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_296 = count >= 10'h1 & count <= _T_27 ? _GEN_196 : L0Memory_67; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_297 = count >= 10'h1 & count <= _T_27 ? _GEN_197 : L0Memory_68; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_298 = count >= 10'h1 & count <= _T_27 ? _GEN_198 : L0Memory_69; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_299 = count >= 10'h1 & count <= _T_27 ? _GEN_199 : L0Memory_70; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_300 = count >= 10'h1 & count <= _T_27 ? _GEN_200 : L0Memory_71; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_301 = count >= 10'h1 & count <= _T_27 ? _GEN_201 : L0Memory_72; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_302 = count >= 10'h1 & count <= _T_27 ? _GEN_202 : L0Memory_73; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_303 = count >= 10'h1 & count <= _T_27 ? _GEN_203 : L0Memory_74; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_304 = count >= 10'h1 & count <= _T_27 ? _GEN_204 : L0Memory_75; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_305 = count >= 10'h1 & count <= _T_27 ? _GEN_205 : L0Memory_76; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_306 = count >= 10'h1 & count <= _T_27 ? _GEN_206 : L0Memory_77; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_307 = count >= 10'h1 & count <= _T_27 ? _GEN_207 : L0Memory_78; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_308 = count >= 10'h1 & count <= _T_27 ? _GEN_208 : L0Memory_79; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_309 = count >= 10'h1 & count <= _T_27 ? _GEN_209 : L0Memory_80; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_310 = count >= 10'h1 & count <= _T_27 ? _GEN_210 : L0Memory_81; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_311 = count >= 10'h1 & count <= _T_27 ? _GEN_211 : L0Memory_82; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_312 = count >= 10'h1 & count <= _T_27 ? _GEN_212 : L0Memory_83; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_313 = count >= 10'h1 & count <= _T_27 ? _GEN_213 : L0Memory_84; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_314 = count >= 10'h1 & count <= _T_27 ? _GEN_214 : L0Memory_85; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_315 = count >= 10'h1 & count <= _T_27 ? _GEN_215 : L0Memory_86; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_316 = count >= 10'h1 & count <= _T_27 ? _GEN_216 : L0Memory_87; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_317 = count >= 10'h1 & count <= _T_27 ? _GEN_217 : L0Memory_88; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_318 = count >= 10'h1 & count <= _T_27 ? _GEN_218 : L0Memory_89; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_319 = count >= 10'h1 & count <= _T_27 ? _GEN_219 : L0Memory_90; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_320 = count >= 10'h1 & count <= _T_27 ? _GEN_220 : L0Memory_91; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_321 = count >= 10'h1 & count <= _T_27 ? _GEN_221 : L0Memory_92; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_322 = count >= 10'h1 & count <= _T_27 ? _GEN_222 : L0Memory_93; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_323 = count >= 10'h1 & count <= _T_27 ? _GEN_223 : L0Memory_94; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_324 = count >= 10'h1 & count <= _T_27 ? _GEN_224 : L0Memory_95; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_325 = count >= 10'h1 & count <= _T_27 ? _GEN_225 : L0Memory_96; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_326 = count >= 10'h1 & count <= _T_27 ? _GEN_226 : L0Memory_97; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_327 = count >= 10'h1 & count <= _T_27 ? _GEN_227 : L0Memory_98; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_328 = count >= 10'h1 & count <= _T_27 ? _GEN_228 : L0Memory_99; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [5:0] _GEN_329 = count >= 10'h1 & count <= _T_27 ? _L0Index_T_2 : _GEN_128; // @[PEArray.scala 198:59 PEArray.scala 200:17]
  wire [9:0] _GEN_330 = count == count_max ? 10'h0 : _GEN_127; // @[PEArray.scala 202:32 PEArray.scala 203:15]
  wire [2:0] _GEN_331 = count == count_max ? 3'h0 : state; // @[PEArray.scala 202:32 PEArray.scala 204:15 PEArray.scala 100:22]
  wire [9:0] _GEN_865 = {{4'd0}, GRU_out_width}; // @[PEArray.scala 220:19]
  wire [9:0] _GEN_0 = count % _GEN_865; // @[PEArray.scala 220:19]
  wire [5:0] _T_36 = _GEN_0[5:0]; // @[PEArray.scala 220:19]
  wire [5:0] _T_38 = GRU_out_width - 6'h1; // @[PEArray.scala 220:55]
  wire [5:0] _GEN_334 = _T_36 == _T_38 ? _L0Index_T_2 : L0index_begin; // @[PEArray.scala 220:62 PEArray.scala 221:17 PEArray.scala 214:15]
  wire [5:0] _GEN_346 = _T_41 ? _GEN_334 : L0Index; // @[Conditional.scala 39:67 PEArray.scala 39:24]
  wire [9:0] _GEN_347 = _T_41 ? _GEN_330 : count; // @[Conditional.scala 39:67 PEArray.scala 101:22]
  wire [2:0] _GEN_348 = _T_41 ? _GEN_331 : state; // @[Conditional.scala 39:67 PEArray.scala 100:22]
  wire [5:0] _GEN_353 = _T_31 ? _GEN_334 : _GEN_346; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_354 = _T_31 ? _GEN_330 : _GEN_347; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_355 = _T_31 ? _GEN_331 : _GEN_348; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_356 = _T_22 ? _GEN_330 : _GEN_354; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_357 = _T_22 ? _GEN_329 : _GEN_353; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_458 = _T_22 ? _GEN_331 : _GEN_355; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_690 = _T_3 ? _GEN_118 : {{2'd0}, GRU_out_width}; // @[Conditional.scala 40:58 PEArray.scala 104:26]
  FP16MulAdder FP16MAC ( // @[PEArray.scala 72:23]
    .io_a(FP16MAC_io_a),
    .io_b(FP16MAC_io_b),
    .io_c(FP16MAC_io_c),
    .io_out(FP16MAC_io_out)
  );
  assign io_ToRightPE = mux3out_reg; // @[PEArray.scala 95:16]
  assign io_ToBelowPE = mux2out_reg; // @[PEArray.scala 94:16]
  assign FP16MAC_io_a = sel1 ? io_FromL1 : io_FromLeftPE; // @[PEArray.scala 50:14 PEArray.scala 50:23 PEArray.scala 51:24]
  assign FP16MAC_io_b = sel5 ? mux4out : _GEN_105; // @[PEArray.scala 77:13 PEArray.scala 78:18 PEArray.scala 81:18]
  assign FP16MAC_io_c = sel5 ? _GEN_105 : mux4out; // @[PEArray.scala 77:13 PEArray.scala 79:18 PEArray.scala 82:18]
  always @(posedge clock) begin
    if (reset) begin // @[PEArray.scala 39:24]
      L0Index <= 6'h0; // @[PEArray.scala 39:24]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h2; // @[PEArray.scala 159:15]
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        L0Index <= 6'hb; // @[PEArray.scala 181:15]
      end else begin
        L0Index <= _GEN_357;
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_0 <= _GEN_229;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_1 <= _GEN_230;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_2 <= _GEN_231;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_3 <= _GEN_232;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_4 <= _GEN_233;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_5 <= _GEN_234;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_6 <= _GEN_235;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_7 <= _GEN_236;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_8 <= _GEN_237;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_9 <= _GEN_238;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_10 <= _GEN_239;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_11 <= _GEN_240;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_12 <= _GEN_241;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_13 <= _GEN_242;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_14 <= _GEN_243;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_15 <= _GEN_244;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_16 <= _GEN_245;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_17 <= _GEN_246;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_18 <= _GEN_247;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_19 <= _GEN_248;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_20 <= _GEN_249;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_21 <= _GEN_250;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_22 <= _GEN_251;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_23 <= _GEN_252;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_24 <= _GEN_253;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_25 <= _GEN_254;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_26 <= _GEN_255;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_27 <= _GEN_256;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_28 <= _GEN_257;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_29 <= _GEN_258;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_30 <= _GEN_259;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_31 <= _GEN_260;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_32 <= _GEN_261;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_33 <= _GEN_262;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_34 <= _GEN_263;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_35 <= _GEN_264;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_36 <= _GEN_265;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_37 <= _GEN_266;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_38 <= _GEN_267;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_39 <= _GEN_268;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_40 <= _GEN_269;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_41 <= _GEN_270;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_42 <= _GEN_271;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_43 <= _GEN_272;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_44 <= _GEN_273;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_45 <= _GEN_274;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_46 <= _GEN_275;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_47 <= _GEN_276;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_48 <= _GEN_277;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_49 <= _GEN_278;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_50 <= _GEN_279;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_51 <= _GEN_280;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_52 <= _GEN_281;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_53 <= _GEN_282;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_54 <= _GEN_283;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_55 <= _GEN_284;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_56 <= _GEN_285;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_57 <= _GEN_286;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_58 <= _GEN_287;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_59 <= _GEN_288;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_60 <= _GEN_289;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_61 <= _GEN_290;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_62 <= _GEN_291;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_63 <= _GEN_292;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_64 <= _GEN_293;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_65 <= _GEN_294;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_66 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_67 <= _GEN_296;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_68 <= _GEN_297;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_69 <= _GEN_298;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_70 <= _GEN_299;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_71 <= _GEN_300;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_72 <= _GEN_301;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_73 <= _GEN_302;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_74 <= _GEN_303;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_75 <= _GEN_304;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_76 <= _GEN_305;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_77 <= _GEN_306;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_78 <= _GEN_307;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_79 <= _GEN_308;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_80 <= _GEN_309;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_81 <= _GEN_310;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_82 <= _GEN_311;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_83 <= _GEN_312;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_84 <= _GEN_313;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_85 <= _GEN_314;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_86 <= _GEN_315;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_87 <= _GEN_316;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_88 <= _GEN_317;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_89 <= _GEN_318;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_90 <= _GEN_319;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_91 <= _GEN_320;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_92 <= _GEN_321;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_93 <= _GEN_322;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_94 <= _GEN_323;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_95 <= _GEN_324;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_96 <= _GEN_325;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_97 <= _GEN_326;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_98 <= _GEN_327;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_99 <= _GEN_328;
          end
        end
      end
    end
    if (reset) begin // @[PEArray.scala 100:22]
      state <= 3'h0; // @[PEArray.scala 100:22]
    end else if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[3]) begin // @[PEArray.scala 116:57]
        if (_T_6) begin // @[Conditional.scala 40:58]
          state <= 3'h0; // @[PEArray.scala 120:19]
        end else begin
          state <= _GEN_113;
        end
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      if (count == 10'h33) begin // @[PEArray.scala 164:27]
        state <= 3'h0; // @[PEArray.scala 166:15]
      end
    end else if (_T_16) begin // @[Conditional.scala 39:67]
      state <= _GEN_126;
    end else begin
      state <= _GEN_458;
    end
    if (reset) begin // @[PEArray.scala 90:28]
      mux2out_reg <= 16'h0; // @[PEArray.scala 90:28]
    end else begin
      mux2out_reg <= MAC_out; // @[PEArray.scala 90:28]
    end
    if (reset) begin // @[PEArray.scala 91:28]
      mux3out_reg <= 16'h0; // @[PEArray.scala 91:28]
    end else if (sel3) begin // @[PEArray.scala 56:14]
      mux3out_reg <= MAC_out; // @[PEArray.scala 56:23]
    end else if (sel1) begin // @[PEArray.scala 50:14]
      mux3out_reg <= io_FromL1; // @[PEArray.scala 50:23]
    end else begin
      mux3out_reg <= io_FromLeftPE; // @[PEArray.scala 51:24]
    end
    if (reset) begin // @[PEArray.scala 101:22]
      count <= 10'h0; // @[PEArray.scala 101:22]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        if (count == 10'h33) begin // @[PEArray.scala 164:27]
          count <= 10'h0; // @[PEArray.scala 165:15]
        end else begin
          count <= _GEN_120;
        end
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        count <= _GEN_125;
      end else begin
        count <= _GEN_356;
      end
    end
    if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[3]) begin // @[PEArray.scala 116:57]
        count_max <= io_control_signal_count; // @[PEArray.scala 143:19]
      end
    end
    if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[3]) begin // @[PEArray.scala 116:57]
        L0index_begin <= io_control_signal_L0index; // @[PEArray.scala 144:23]
      end
    end
    GRU_out_width <= _GEN_690[5:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  L0Index = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  L0Memory_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  L0Memory_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  L0Memory_2 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  L0Memory_3 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  L0Memory_4 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  L0Memory_5 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  L0Memory_6 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  L0Memory_7 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  L0Memory_8 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  L0Memory_9 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  L0Memory_10 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  L0Memory_11 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  L0Memory_12 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  L0Memory_13 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  L0Memory_14 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  L0Memory_15 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  L0Memory_16 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  L0Memory_17 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  L0Memory_18 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  L0Memory_19 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  L0Memory_20 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  L0Memory_21 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  L0Memory_22 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  L0Memory_23 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  L0Memory_24 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  L0Memory_25 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  L0Memory_26 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  L0Memory_27 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  L0Memory_28 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  L0Memory_29 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  L0Memory_30 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  L0Memory_31 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  L0Memory_32 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  L0Memory_33 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  L0Memory_34 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  L0Memory_35 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  L0Memory_36 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  L0Memory_37 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  L0Memory_38 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  L0Memory_39 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  L0Memory_40 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  L0Memory_41 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  L0Memory_42 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  L0Memory_43 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  L0Memory_44 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  L0Memory_45 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  L0Memory_46 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  L0Memory_47 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  L0Memory_48 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  L0Memory_49 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  L0Memory_50 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  L0Memory_51 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  L0Memory_52 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  L0Memory_53 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  L0Memory_54 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  L0Memory_55 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  L0Memory_56 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  L0Memory_57 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  L0Memory_58 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  L0Memory_59 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  L0Memory_60 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  L0Memory_61 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  L0Memory_62 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  L0Memory_63 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  L0Memory_64 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  L0Memory_65 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  L0Memory_66 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  L0Memory_67 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  L0Memory_68 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  L0Memory_69 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  L0Memory_70 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  L0Memory_71 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  L0Memory_72 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  L0Memory_73 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  L0Memory_74 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  L0Memory_75 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  L0Memory_76 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  L0Memory_77 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  L0Memory_78 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  L0Memory_79 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  L0Memory_80 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  L0Memory_81 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  L0Memory_82 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  L0Memory_83 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  L0Memory_84 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  L0Memory_85 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  L0Memory_86 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  L0Memory_87 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  L0Memory_88 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  L0Memory_89 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  L0Memory_90 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  L0Memory_91 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  L0Memory_92 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  L0Memory_93 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  L0Memory_94 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  L0Memory_95 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  L0Memory_96 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  L0Memory_97 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  L0Memory_98 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  L0Memory_99 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  state = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  mux2out_reg = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  mux3out_reg = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  count = _RAND_104[9:0];
  _RAND_105 = {1{`RANDOM}};
  count_max = _RAND_105[9:0];
  _RAND_106 = {1{`RANDOM}};
  L0index_begin = _RAND_106[5:0];
  _RAND_107 = {1{`RANDOM}};
  GRU_out_width = _RAND_107[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PE_27(
  input         clock,
  input         reset,
  input  [15:0] io_FromAbovePE,
  input  [15:0] io_FromLeftPE,
  input  [15:0] io_FromL1,
  input  [11:0] io_control_signal_mask,
  output [15:0] io_ToRightPE,
  output [15:0] io_ToBelowPE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] FP16MAC_io_a; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_b; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_c; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_out; // @[PEArray.scala 72:23]
  reg [5:0] L0Index; // @[PEArray.scala 39:24]
  reg [15:0] L0Memory_0; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_1; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_2; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_3; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_4; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_5; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_6; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_7; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_8; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_9; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_10; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_11; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_12; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_13; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_14; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_15; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_16; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_17; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_18; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_19; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_20; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_21; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_22; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_23; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_24; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_25; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_26; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_27; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_28; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_29; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_30; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_31; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_32; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_33; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_34; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_35; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_36; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_37; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_38; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_39; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_40; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_41; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_42; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_43; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_44; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_45; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_46; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_47; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_48; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_49; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_50; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_51; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_52; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_53; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_54; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_55; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_56; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_57; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_58; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_59; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_60; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_61; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_62; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_63; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_64; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_65; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_66; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_67; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_68; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_69; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_70; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_71; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_72; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_73; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_74; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_75; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_76; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_77; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_78; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_79; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_80; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_81; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_82; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_83; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_84; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_85; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_86; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_87; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_88; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_89; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_90; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_91; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_92; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_93; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_94; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_95; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_96; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_97; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_98; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_99; // @[PEArray.scala 40:21]
  reg [2:0] state; // @[PEArray.scala 100:22]
  wire  _T_3 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_12 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_16 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_22 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_31 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_41 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_342 = _T_41 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 231:12 PEArray.scala 32:8]
  wire  _GEN_349 = _T_31 ? 1'h0 : _GEN_342; // @[Conditional.scala 39:67 PEArray.scala 208:12]
  wire  _GEN_459 = _T_22 | _GEN_349; // @[Conditional.scala 39:67 PEArray.scala 32:8]
  wire  _GEN_463 = _T_16 ? 1'h0 : _GEN_459; // @[Conditional.scala 39:67]
  wire  _GEN_572 = _T_12 | _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 149:12]
  wire  sel1 = _T_3 | _GEN_572; // @[Conditional.scala 40:58 PEArray.scala 108:12]
  wire [15:0] MAC_out = FP16MAC_io_out; // @[PEArray.scala 47:21 PEArray.scala 85:11]
  wire  _GEN_465 = _T_16 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 177:12]
  wire  _GEN_580 = _T_12 | _GEN_465; // @[Conditional.scala 39:67 PEArray.scala 34:8]
  wire  sel3 = _T_3 | _GEN_580; // @[Conditional.scala 40:58 PEArray.scala 110:12]
  wire [1:0] _GEN_344 = _T_41 ? 2'h2 : 2'h0; // @[Conditional.scala 39:67 PEArray.scala 233:12 PEArray.scala 35:8]
  wire [1:0] _GEN_351 = _T_31 ? 2'h2 : _GEN_344; // @[Conditional.scala 39:67 PEArray.scala 210:12]
  wire [1:0] _GEN_461 = _T_22 ? 2'h0 : _GEN_351; // @[Conditional.scala 39:67 PEArray.scala 35:8]
  wire [1:0] _GEN_466 = _T_16 ? 2'h0 : _GEN_461; // @[Conditional.scala 39:67 PEArray.scala 178:12]
  wire [1:0] _GEN_574 = _T_12 ? 2'h0 : _GEN_466; // @[Conditional.scala 39:67]
  wire [1:0] sel4 = _T_3 ? 2'h0 : _GEN_574; // @[Conditional.scala 40:58 PEArray.scala 111:12]
  wire [15:0] _GEN_3 = sel4 == 2'h2 ? io_FromL1 : 16'h0; // @[PEArray.scala 65:28 PEArray.scala 66:15 PEArray.scala 69:15]
  wire [15:0] _GEN_4 = sel4 == 2'h1 ? io_FromAbovePE : _GEN_3; // @[PEArray.scala 62:28 PEArray.scala 63:15]
  wire [15:0] mux4out = sel4 == 2'h0 ? 16'h0 : _GEN_4; // @[PEArray.scala 59:22 PEArray.scala 60:13]
  wire [15:0] _GEN_7 = 6'h1 == L0Index ? L0Memory_1 : L0Memory_0; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_8 = 6'h2 == L0Index ? L0Memory_2 : _GEN_7; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_9 = 6'h3 == L0Index ? L0Memory_3 : _GEN_8; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_10 = 6'h4 == L0Index ? L0Memory_4 : _GEN_9; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_11 = 6'h5 == L0Index ? L0Memory_5 : _GEN_10; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_12 = 6'h6 == L0Index ? L0Memory_6 : _GEN_11; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_13 = 6'h7 == L0Index ? L0Memory_7 : _GEN_12; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_14 = 6'h8 == L0Index ? L0Memory_8 : _GEN_13; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_15 = 6'h9 == L0Index ? L0Memory_9 : _GEN_14; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_16 = 6'ha == L0Index ? L0Memory_10 : _GEN_15; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_17 = 6'hb == L0Index ? L0Memory_11 : _GEN_16; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_18 = 6'hc == L0Index ? L0Memory_12 : _GEN_17; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_19 = 6'hd == L0Index ? L0Memory_13 : _GEN_18; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_20 = 6'he == L0Index ? L0Memory_14 : _GEN_19; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_21 = 6'hf == L0Index ? L0Memory_15 : _GEN_20; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_22 = 6'h10 == L0Index ? L0Memory_16 : _GEN_21; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_23 = 6'h11 == L0Index ? L0Memory_17 : _GEN_22; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_24 = 6'h12 == L0Index ? L0Memory_18 : _GEN_23; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_25 = 6'h13 == L0Index ? L0Memory_19 : _GEN_24; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_26 = 6'h14 == L0Index ? L0Memory_20 : _GEN_25; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_27 = 6'h15 == L0Index ? L0Memory_21 : _GEN_26; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_28 = 6'h16 == L0Index ? L0Memory_22 : _GEN_27; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_29 = 6'h17 == L0Index ? L0Memory_23 : _GEN_28; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_30 = 6'h18 == L0Index ? L0Memory_24 : _GEN_29; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_31 = 6'h19 == L0Index ? L0Memory_25 : _GEN_30; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_32 = 6'h1a == L0Index ? L0Memory_26 : _GEN_31; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_33 = 6'h1b == L0Index ? L0Memory_27 : _GEN_32; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_34 = 6'h1c == L0Index ? L0Memory_28 : _GEN_33; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_35 = 6'h1d == L0Index ? L0Memory_29 : _GEN_34; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_36 = 6'h1e == L0Index ? L0Memory_30 : _GEN_35; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_37 = 6'h1f == L0Index ? L0Memory_31 : _GEN_36; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_38 = 6'h20 == L0Index ? L0Memory_32 : _GEN_37; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_39 = 6'h21 == L0Index ? L0Memory_33 : _GEN_38; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_40 = 6'h22 == L0Index ? L0Memory_34 : _GEN_39; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_41 = 6'h23 == L0Index ? L0Memory_35 : _GEN_40; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_42 = 6'h24 == L0Index ? L0Memory_36 : _GEN_41; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_43 = 6'h25 == L0Index ? L0Memory_37 : _GEN_42; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_44 = 6'h26 == L0Index ? L0Memory_38 : _GEN_43; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_45 = 6'h27 == L0Index ? L0Memory_39 : _GEN_44; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_46 = 6'h28 == L0Index ? L0Memory_40 : _GEN_45; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_47 = 6'h29 == L0Index ? L0Memory_41 : _GEN_46; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_48 = 6'h2a == L0Index ? L0Memory_42 : _GEN_47; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_49 = 6'h2b == L0Index ? L0Memory_43 : _GEN_48; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_50 = 6'h2c == L0Index ? L0Memory_44 : _GEN_49; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_51 = 6'h2d == L0Index ? L0Memory_45 : _GEN_50; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_52 = 6'h2e == L0Index ? L0Memory_46 : _GEN_51; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_53 = 6'h2f == L0Index ? L0Memory_47 : _GEN_52; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_54 = 6'h30 == L0Index ? L0Memory_48 : _GEN_53; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_55 = 6'h31 == L0Index ? L0Memory_49 : _GEN_54; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_56 = 6'h32 == L0Index ? L0Memory_50 : _GEN_55; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_57 = 6'h33 == L0Index ? L0Memory_51 : _GEN_56; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_58 = 6'h34 == L0Index ? L0Memory_52 : _GEN_57; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_59 = 6'h35 == L0Index ? L0Memory_53 : _GEN_58; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_60 = 6'h36 == L0Index ? L0Memory_54 : _GEN_59; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_61 = 6'h37 == L0Index ? L0Memory_55 : _GEN_60; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_62 = 6'h38 == L0Index ? L0Memory_56 : _GEN_61; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_63 = 6'h39 == L0Index ? L0Memory_57 : _GEN_62; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_64 = 6'h3a == L0Index ? L0Memory_58 : _GEN_63; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_65 = 6'h3b == L0Index ? L0Memory_59 : _GEN_64; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_66 = 6'h3c == L0Index ? L0Memory_60 : _GEN_65; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_67 = 6'h3d == L0Index ? L0Memory_61 : _GEN_66; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_68 = 6'h3e == L0Index ? L0Memory_62 : _GEN_67; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_69 = 6'h3f == L0Index ? L0Memory_63 : _GEN_68; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [6:0] _GEN_793 = {{1'd0}, L0Index}; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_70 = 7'h40 == _GEN_793 ? L0Memory_64 : _GEN_69; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_71 = 7'h41 == _GEN_793 ? L0Memory_65 : _GEN_70; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_72 = 7'h42 == _GEN_793 ? L0Memory_66 : _GEN_71; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_73 = 7'h43 == _GEN_793 ? L0Memory_67 : _GEN_72; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_74 = 7'h44 == _GEN_793 ? L0Memory_68 : _GEN_73; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_75 = 7'h45 == _GEN_793 ? L0Memory_69 : _GEN_74; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_76 = 7'h46 == _GEN_793 ? L0Memory_70 : _GEN_75; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_77 = 7'h47 == _GEN_793 ? L0Memory_71 : _GEN_76; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_78 = 7'h48 == _GEN_793 ? L0Memory_72 : _GEN_77; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_79 = 7'h49 == _GEN_793 ? L0Memory_73 : _GEN_78; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_80 = 7'h4a == _GEN_793 ? L0Memory_74 : _GEN_79; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_81 = 7'h4b == _GEN_793 ? L0Memory_75 : _GEN_80; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_82 = 7'h4c == _GEN_793 ? L0Memory_76 : _GEN_81; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_83 = 7'h4d == _GEN_793 ? L0Memory_77 : _GEN_82; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_84 = 7'h4e == _GEN_793 ? L0Memory_78 : _GEN_83; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_85 = 7'h4f == _GEN_793 ? L0Memory_79 : _GEN_84; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_86 = 7'h50 == _GEN_793 ? L0Memory_80 : _GEN_85; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_87 = 7'h51 == _GEN_793 ? L0Memory_81 : _GEN_86; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_88 = 7'h52 == _GEN_793 ? L0Memory_82 : _GEN_87; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_89 = 7'h53 == _GEN_793 ? L0Memory_83 : _GEN_88; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_90 = 7'h54 == _GEN_793 ? L0Memory_84 : _GEN_89; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_91 = 7'h55 == _GEN_793 ? L0Memory_85 : _GEN_90; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_92 = 7'h56 == _GEN_793 ? L0Memory_86 : _GEN_91; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_93 = 7'h57 == _GEN_793 ? L0Memory_87 : _GEN_92; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_94 = 7'h58 == _GEN_793 ? L0Memory_88 : _GEN_93; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_95 = 7'h59 == _GEN_793 ? L0Memory_89 : _GEN_94; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_96 = 7'h5a == _GEN_793 ? L0Memory_90 : _GEN_95; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_97 = 7'h5b == _GEN_793 ? L0Memory_91 : _GEN_96; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_98 = 7'h5c == _GEN_793 ? L0Memory_92 : _GEN_97; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_99 = 7'h5d == _GEN_793 ? L0Memory_93 : _GEN_98; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_100 = 7'h5e == _GEN_793 ? L0Memory_94 : _GEN_99; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_101 = 7'h5f == _GEN_793 ? L0Memory_95 : _GEN_100; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_102 = 7'h60 == _GEN_793 ? L0Memory_96 : _GEN_101; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_103 = 7'h61 == _GEN_793 ? L0Memory_97 : _GEN_102; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_104 = 7'h62 == _GEN_793 ? L0Memory_98 : _GEN_103; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_105 = 7'h63 == _GEN_793 ? L0Memory_99 : _GEN_104; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire  _GEN_575 = _T_12 ? 1'h0 : _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 157:12]
  wire  sel5 = _T_3 ? 1'h0 : _GEN_575; // @[Conditional.scala 40:58 PEArray.scala 112:12]
  reg [15:0] mux2out_reg; // @[PEArray.scala 90:28]
  reg [15:0] mux3out_reg; // @[PEArray.scala 91:28]
  reg [9:0] count; // @[PEArray.scala 101:22]
  reg [5:0] GRU_out_width; // @[PEArray.scala 104:26]
  wire [7:0] _GEN_118 = io_control_signal_mask[2] ? 8'h0 : {{2'd0}, GRU_out_width}; // @[PEArray.scala 116:57 PEArray.scala 145:23 PEArray.scala 104:26]
  wire [9:0] _count_T_1 = count + 10'h1; // @[PEArray.scala 162:24]
  wire [9:0] _GEN_120 = count != 10'h33 ? _count_T_1 : count; // @[PEArray.scala 161:27 PEArray.scala 162:15 PEArray.scala 101:22]
  wire [9:0] _GEN_124 = count != 10'h188 ? _count_T_1 : count; // @[PEArray.scala 183:28 PEArray.scala 184:15 PEArray.scala 101:22]
  wire [9:0] _GEN_125 = count == 10'h188 ? 10'h0 : _GEN_124; // @[PEArray.scala 186:28 PEArray.scala 187:15]
  wire [2:0] _GEN_126 = count == 10'h188 ? 3'h0 : state; // @[PEArray.scala 186:28 PEArray.scala 188:15 PEArray.scala 100:22]
  wire [9:0] _GEN_127 = count != 10'h0 ? _count_T_1 : count; // @[PEArray.scala 192:32 PEArray.scala 193:15 PEArray.scala 101:22]
  wire  _T_24 = count == 10'h0; // @[PEArray.scala 195:18]
  wire [5:0] _GEN_128 = count == 10'h0 ? 6'h0 : L0Index; // @[PEArray.scala 195:26 PEArray.scala 196:17 PEArray.scala 39:24]
  wire [9:0] _T_27 = 10'h0 - 10'h1; // @[PEArray.scala 198:51]
  wire [15:0] _GEN_129 = 6'h0 == L0Index ? io_FromL1 : L0Memory_0; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_130 = 6'h1 == L0Index ? io_FromL1 : L0Memory_1; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_131 = 6'h2 == L0Index ? io_FromL1 : L0Memory_2; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_132 = 6'h3 == L0Index ? io_FromL1 : L0Memory_3; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_133 = 6'h4 == L0Index ? io_FromL1 : L0Memory_4; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_134 = 6'h5 == L0Index ? io_FromL1 : L0Memory_5; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_135 = 6'h6 == L0Index ? io_FromL1 : L0Memory_6; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_136 = 6'h7 == L0Index ? io_FromL1 : L0Memory_7; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_137 = 6'h8 == L0Index ? io_FromL1 : L0Memory_8; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_138 = 6'h9 == L0Index ? io_FromL1 : L0Memory_9; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_139 = 6'ha == L0Index ? io_FromL1 : L0Memory_10; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_140 = 6'hb == L0Index ? io_FromL1 : L0Memory_11; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_141 = 6'hc == L0Index ? io_FromL1 : L0Memory_12; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_142 = 6'hd == L0Index ? io_FromL1 : L0Memory_13; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_143 = 6'he == L0Index ? io_FromL1 : L0Memory_14; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_144 = 6'hf == L0Index ? io_FromL1 : L0Memory_15; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_145 = 6'h10 == L0Index ? io_FromL1 : L0Memory_16; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_146 = 6'h11 == L0Index ? io_FromL1 : L0Memory_17; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_147 = 6'h12 == L0Index ? io_FromL1 : L0Memory_18; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_148 = 6'h13 == L0Index ? io_FromL1 : L0Memory_19; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_149 = 6'h14 == L0Index ? io_FromL1 : L0Memory_20; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_150 = 6'h15 == L0Index ? io_FromL1 : L0Memory_21; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_151 = 6'h16 == L0Index ? io_FromL1 : L0Memory_22; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_152 = 6'h17 == L0Index ? io_FromL1 : L0Memory_23; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_153 = 6'h18 == L0Index ? io_FromL1 : L0Memory_24; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_154 = 6'h19 == L0Index ? io_FromL1 : L0Memory_25; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_155 = 6'h1a == L0Index ? io_FromL1 : L0Memory_26; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_156 = 6'h1b == L0Index ? io_FromL1 : L0Memory_27; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_157 = 6'h1c == L0Index ? io_FromL1 : L0Memory_28; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_158 = 6'h1d == L0Index ? io_FromL1 : L0Memory_29; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_159 = 6'h1e == L0Index ? io_FromL1 : L0Memory_30; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_160 = 6'h1f == L0Index ? io_FromL1 : L0Memory_31; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_161 = 6'h20 == L0Index ? io_FromL1 : L0Memory_32; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_162 = 6'h21 == L0Index ? io_FromL1 : L0Memory_33; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_163 = 6'h22 == L0Index ? io_FromL1 : L0Memory_34; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_164 = 6'h23 == L0Index ? io_FromL1 : L0Memory_35; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_165 = 6'h24 == L0Index ? io_FromL1 : L0Memory_36; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_166 = 6'h25 == L0Index ? io_FromL1 : L0Memory_37; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_167 = 6'h26 == L0Index ? io_FromL1 : L0Memory_38; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_168 = 6'h27 == L0Index ? io_FromL1 : L0Memory_39; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_169 = 6'h28 == L0Index ? io_FromL1 : L0Memory_40; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_170 = 6'h29 == L0Index ? io_FromL1 : L0Memory_41; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_171 = 6'h2a == L0Index ? io_FromL1 : L0Memory_42; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_172 = 6'h2b == L0Index ? io_FromL1 : L0Memory_43; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_173 = 6'h2c == L0Index ? io_FromL1 : L0Memory_44; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_174 = 6'h2d == L0Index ? io_FromL1 : L0Memory_45; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_175 = 6'h2e == L0Index ? io_FromL1 : L0Memory_46; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_176 = 6'h2f == L0Index ? io_FromL1 : L0Memory_47; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_177 = 6'h30 == L0Index ? io_FromL1 : L0Memory_48; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_178 = 6'h31 == L0Index ? io_FromL1 : L0Memory_49; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_179 = 6'h32 == L0Index ? io_FromL1 : L0Memory_50; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_180 = 6'h33 == L0Index ? io_FromL1 : L0Memory_51; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_181 = 6'h34 == L0Index ? io_FromL1 : L0Memory_52; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_182 = 6'h35 == L0Index ? io_FromL1 : L0Memory_53; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_183 = 6'h36 == L0Index ? io_FromL1 : L0Memory_54; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_184 = 6'h37 == L0Index ? io_FromL1 : L0Memory_55; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_185 = 6'h38 == L0Index ? io_FromL1 : L0Memory_56; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_186 = 6'h39 == L0Index ? io_FromL1 : L0Memory_57; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_187 = 6'h3a == L0Index ? io_FromL1 : L0Memory_58; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_188 = 6'h3b == L0Index ? io_FromL1 : L0Memory_59; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_189 = 6'h3c == L0Index ? io_FromL1 : L0Memory_60; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_190 = 6'h3d == L0Index ? io_FromL1 : L0Memory_61; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_191 = 6'h3e == L0Index ? io_FromL1 : L0Memory_62; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_192 = 6'h3f == L0Index ? io_FromL1 : L0Memory_63; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_193 = 7'h40 == _GEN_793 ? io_FromL1 : L0Memory_64; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_194 = 7'h41 == _GEN_793 ? io_FromL1 : L0Memory_65; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_195 = 7'h42 == _GEN_793 ? io_FromL1 : L0Memory_66; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_196 = 7'h43 == _GEN_793 ? io_FromL1 : L0Memory_67; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_197 = 7'h44 == _GEN_793 ? io_FromL1 : L0Memory_68; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_198 = 7'h45 == _GEN_793 ? io_FromL1 : L0Memory_69; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_199 = 7'h46 == _GEN_793 ? io_FromL1 : L0Memory_70; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_200 = 7'h47 == _GEN_793 ? io_FromL1 : L0Memory_71; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_201 = 7'h48 == _GEN_793 ? io_FromL1 : L0Memory_72; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_202 = 7'h49 == _GEN_793 ? io_FromL1 : L0Memory_73; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_203 = 7'h4a == _GEN_793 ? io_FromL1 : L0Memory_74; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_204 = 7'h4b == _GEN_793 ? io_FromL1 : L0Memory_75; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_205 = 7'h4c == _GEN_793 ? io_FromL1 : L0Memory_76; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_206 = 7'h4d == _GEN_793 ? io_FromL1 : L0Memory_77; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_207 = 7'h4e == _GEN_793 ? io_FromL1 : L0Memory_78; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_208 = 7'h4f == _GEN_793 ? io_FromL1 : L0Memory_79; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_209 = 7'h50 == _GEN_793 ? io_FromL1 : L0Memory_80; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_210 = 7'h51 == _GEN_793 ? io_FromL1 : L0Memory_81; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_211 = 7'h52 == _GEN_793 ? io_FromL1 : L0Memory_82; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_212 = 7'h53 == _GEN_793 ? io_FromL1 : L0Memory_83; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_213 = 7'h54 == _GEN_793 ? io_FromL1 : L0Memory_84; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_214 = 7'h55 == _GEN_793 ? io_FromL1 : L0Memory_85; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_215 = 7'h56 == _GEN_793 ? io_FromL1 : L0Memory_86; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_216 = 7'h57 == _GEN_793 ? io_FromL1 : L0Memory_87; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_217 = 7'h58 == _GEN_793 ? io_FromL1 : L0Memory_88; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_218 = 7'h59 == _GEN_793 ? io_FromL1 : L0Memory_89; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_219 = 7'h5a == _GEN_793 ? io_FromL1 : L0Memory_90; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_220 = 7'h5b == _GEN_793 ? io_FromL1 : L0Memory_91; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_221 = 7'h5c == _GEN_793 ? io_FromL1 : L0Memory_92; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_222 = 7'h5d == _GEN_793 ? io_FromL1 : L0Memory_93; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_223 = 7'h5e == _GEN_793 ? io_FromL1 : L0Memory_94; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_224 = 7'h5f == _GEN_793 ? io_FromL1 : L0Memory_95; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_225 = 7'h60 == _GEN_793 ? io_FromL1 : L0Memory_96; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_226 = 7'h61 == _GEN_793 ? io_FromL1 : L0Memory_97; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_227 = 7'h62 == _GEN_793 ? io_FromL1 : L0Memory_98; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_228 = 7'h63 == _GEN_793 ? io_FromL1 : L0Memory_99; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [5:0] _L0Index_T_2 = L0Index + 6'h1; // @[PEArray.scala 200:28]
  wire [15:0] _GEN_229 = count >= 10'h1 & count <= _T_27 ? _GEN_129 : L0Memory_0; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_230 = count >= 10'h1 & count <= _T_27 ? _GEN_130 : L0Memory_1; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_231 = count >= 10'h1 & count <= _T_27 ? _GEN_131 : L0Memory_2; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_232 = count >= 10'h1 & count <= _T_27 ? _GEN_132 : L0Memory_3; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_233 = count >= 10'h1 & count <= _T_27 ? _GEN_133 : L0Memory_4; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_234 = count >= 10'h1 & count <= _T_27 ? _GEN_134 : L0Memory_5; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_235 = count >= 10'h1 & count <= _T_27 ? _GEN_135 : L0Memory_6; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_236 = count >= 10'h1 & count <= _T_27 ? _GEN_136 : L0Memory_7; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_237 = count >= 10'h1 & count <= _T_27 ? _GEN_137 : L0Memory_8; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_238 = count >= 10'h1 & count <= _T_27 ? _GEN_138 : L0Memory_9; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_239 = count >= 10'h1 & count <= _T_27 ? _GEN_139 : L0Memory_10; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_240 = count >= 10'h1 & count <= _T_27 ? _GEN_140 : L0Memory_11; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_241 = count >= 10'h1 & count <= _T_27 ? _GEN_141 : L0Memory_12; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_242 = count >= 10'h1 & count <= _T_27 ? _GEN_142 : L0Memory_13; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_243 = count >= 10'h1 & count <= _T_27 ? _GEN_143 : L0Memory_14; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_244 = count >= 10'h1 & count <= _T_27 ? _GEN_144 : L0Memory_15; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_245 = count >= 10'h1 & count <= _T_27 ? _GEN_145 : L0Memory_16; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_246 = count >= 10'h1 & count <= _T_27 ? _GEN_146 : L0Memory_17; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_247 = count >= 10'h1 & count <= _T_27 ? _GEN_147 : L0Memory_18; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_248 = count >= 10'h1 & count <= _T_27 ? _GEN_148 : L0Memory_19; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_249 = count >= 10'h1 & count <= _T_27 ? _GEN_149 : L0Memory_20; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_250 = count >= 10'h1 & count <= _T_27 ? _GEN_150 : L0Memory_21; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_251 = count >= 10'h1 & count <= _T_27 ? _GEN_151 : L0Memory_22; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_252 = count >= 10'h1 & count <= _T_27 ? _GEN_152 : L0Memory_23; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_253 = count >= 10'h1 & count <= _T_27 ? _GEN_153 : L0Memory_24; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_254 = count >= 10'h1 & count <= _T_27 ? _GEN_154 : L0Memory_25; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_255 = count >= 10'h1 & count <= _T_27 ? _GEN_155 : L0Memory_26; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_256 = count >= 10'h1 & count <= _T_27 ? _GEN_156 : L0Memory_27; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_257 = count >= 10'h1 & count <= _T_27 ? _GEN_157 : L0Memory_28; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_258 = count >= 10'h1 & count <= _T_27 ? _GEN_158 : L0Memory_29; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_259 = count >= 10'h1 & count <= _T_27 ? _GEN_159 : L0Memory_30; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_260 = count >= 10'h1 & count <= _T_27 ? _GEN_160 : L0Memory_31; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_261 = count >= 10'h1 & count <= _T_27 ? _GEN_161 : L0Memory_32; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_262 = count >= 10'h1 & count <= _T_27 ? _GEN_162 : L0Memory_33; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_263 = count >= 10'h1 & count <= _T_27 ? _GEN_163 : L0Memory_34; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_264 = count >= 10'h1 & count <= _T_27 ? _GEN_164 : L0Memory_35; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_265 = count >= 10'h1 & count <= _T_27 ? _GEN_165 : L0Memory_36; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_266 = count >= 10'h1 & count <= _T_27 ? _GEN_166 : L0Memory_37; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_267 = count >= 10'h1 & count <= _T_27 ? _GEN_167 : L0Memory_38; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_268 = count >= 10'h1 & count <= _T_27 ? _GEN_168 : L0Memory_39; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_269 = count >= 10'h1 & count <= _T_27 ? _GEN_169 : L0Memory_40; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_270 = count >= 10'h1 & count <= _T_27 ? _GEN_170 : L0Memory_41; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_271 = count >= 10'h1 & count <= _T_27 ? _GEN_171 : L0Memory_42; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_272 = count >= 10'h1 & count <= _T_27 ? _GEN_172 : L0Memory_43; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_273 = count >= 10'h1 & count <= _T_27 ? _GEN_173 : L0Memory_44; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_274 = count >= 10'h1 & count <= _T_27 ? _GEN_174 : L0Memory_45; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_275 = count >= 10'h1 & count <= _T_27 ? _GEN_175 : L0Memory_46; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_276 = count >= 10'h1 & count <= _T_27 ? _GEN_176 : L0Memory_47; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_277 = count >= 10'h1 & count <= _T_27 ? _GEN_177 : L0Memory_48; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_278 = count >= 10'h1 & count <= _T_27 ? _GEN_178 : L0Memory_49; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_279 = count >= 10'h1 & count <= _T_27 ? _GEN_179 : L0Memory_50; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_280 = count >= 10'h1 & count <= _T_27 ? _GEN_180 : L0Memory_51; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_281 = count >= 10'h1 & count <= _T_27 ? _GEN_181 : L0Memory_52; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_282 = count >= 10'h1 & count <= _T_27 ? _GEN_182 : L0Memory_53; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_283 = count >= 10'h1 & count <= _T_27 ? _GEN_183 : L0Memory_54; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_284 = count >= 10'h1 & count <= _T_27 ? _GEN_184 : L0Memory_55; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_285 = count >= 10'h1 & count <= _T_27 ? _GEN_185 : L0Memory_56; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_286 = count >= 10'h1 & count <= _T_27 ? _GEN_186 : L0Memory_57; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_287 = count >= 10'h1 & count <= _T_27 ? _GEN_187 : L0Memory_58; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_288 = count >= 10'h1 & count <= _T_27 ? _GEN_188 : L0Memory_59; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_289 = count >= 10'h1 & count <= _T_27 ? _GEN_189 : L0Memory_60; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_290 = count >= 10'h1 & count <= _T_27 ? _GEN_190 : L0Memory_61; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_291 = count >= 10'h1 & count <= _T_27 ? _GEN_191 : L0Memory_62; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_292 = count >= 10'h1 & count <= _T_27 ? _GEN_192 : L0Memory_63; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_293 = count >= 10'h1 & count <= _T_27 ? _GEN_193 : L0Memory_64; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_294 = count >= 10'h1 & count <= _T_27 ? _GEN_194 : L0Memory_65; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_295 = count >= 10'h1 & count <= _T_27 ? _GEN_195 : L0Memory_66; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_296 = count >= 10'h1 & count <= _T_27 ? _GEN_196 : L0Memory_67; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_297 = count >= 10'h1 & count <= _T_27 ? _GEN_197 : L0Memory_68; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_298 = count >= 10'h1 & count <= _T_27 ? _GEN_198 : L0Memory_69; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_299 = count >= 10'h1 & count <= _T_27 ? _GEN_199 : L0Memory_70; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_300 = count >= 10'h1 & count <= _T_27 ? _GEN_200 : L0Memory_71; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_301 = count >= 10'h1 & count <= _T_27 ? _GEN_201 : L0Memory_72; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_302 = count >= 10'h1 & count <= _T_27 ? _GEN_202 : L0Memory_73; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_303 = count >= 10'h1 & count <= _T_27 ? _GEN_203 : L0Memory_74; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_304 = count >= 10'h1 & count <= _T_27 ? _GEN_204 : L0Memory_75; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_305 = count >= 10'h1 & count <= _T_27 ? _GEN_205 : L0Memory_76; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_306 = count >= 10'h1 & count <= _T_27 ? _GEN_206 : L0Memory_77; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_307 = count >= 10'h1 & count <= _T_27 ? _GEN_207 : L0Memory_78; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_308 = count >= 10'h1 & count <= _T_27 ? _GEN_208 : L0Memory_79; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_309 = count >= 10'h1 & count <= _T_27 ? _GEN_209 : L0Memory_80; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_310 = count >= 10'h1 & count <= _T_27 ? _GEN_210 : L0Memory_81; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_311 = count >= 10'h1 & count <= _T_27 ? _GEN_211 : L0Memory_82; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_312 = count >= 10'h1 & count <= _T_27 ? _GEN_212 : L0Memory_83; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_313 = count >= 10'h1 & count <= _T_27 ? _GEN_213 : L0Memory_84; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_314 = count >= 10'h1 & count <= _T_27 ? _GEN_214 : L0Memory_85; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_315 = count >= 10'h1 & count <= _T_27 ? _GEN_215 : L0Memory_86; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_316 = count >= 10'h1 & count <= _T_27 ? _GEN_216 : L0Memory_87; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_317 = count >= 10'h1 & count <= _T_27 ? _GEN_217 : L0Memory_88; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_318 = count >= 10'h1 & count <= _T_27 ? _GEN_218 : L0Memory_89; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_319 = count >= 10'h1 & count <= _T_27 ? _GEN_219 : L0Memory_90; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_320 = count >= 10'h1 & count <= _T_27 ? _GEN_220 : L0Memory_91; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_321 = count >= 10'h1 & count <= _T_27 ? _GEN_221 : L0Memory_92; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_322 = count >= 10'h1 & count <= _T_27 ? _GEN_222 : L0Memory_93; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_323 = count >= 10'h1 & count <= _T_27 ? _GEN_223 : L0Memory_94; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_324 = count >= 10'h1 & count <= _T_27 ? _GEN_224 : L0Memory_95; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_325 = count >= 10'h1 & count <= _T_27 ? _GEN_225 : L0Memory_96; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_326 = count >= 10'h1 & count <= _T_27 ? _GEN_226 : L0Memory_97; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_327 = count >= 10'h1 & count <= _T_27 ? _GEN_227 : L0Memory_98; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_328 = count >= 10'h1 & count <= _T_27 ? _GEN_228 : L0Memory_99; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [5:0] _GEN_329 = count >= 10'h1 & count <= _T_27 ? _L0Index_T_2 : _GEN_128; // @[PEArray.scala 198:59 PEArray.scala 200:17]
  wire [9:0] _GEN_330 = _T_24 ? 10'h0 : _GEN_127; // @[PEArray.scala 202:32 PEArray.scala 203:15]
  wire [2:0] _GEN_331 = _T_24 ? 3'h0 : state; // @[PEArray.scala 202:32 PEArray.scala 204:15 PEArray.scala 100:22]
  wire [9:0] _GEN_865 = {{4'd0}, GRU_out_width}; // @[PEArray.scala 220:19]
  wire [9:0] _GEN_0 = count % _GEN_865; // @[PEArray.scala 220:19]
  wire [5:0] _T_36 = _GEN_0[5:0]; // @[PEArray.scala 220:19]
  wire [5:0] _T_38 = GRU_out_width - 6'h1; // @[PEArray.scala 220:55]
  wire [5:0] _GEN_334 = _T_36 == _T_38 ? _L0Index_T_2 : 6'h0; // @[PEArray.scala 220:62 PEArray.scala 221:17 PEArray.scala 214:15]
  wire [5:0] _GEN_346 = _T_41 ? _GEN_334 : L0Index; // @[Conditional.scala 39:67 PEArray.scala 39:24]
  wire [9:0] _GEN_347 = _T_41 ? _GEN_330 : count; // @[Conditional.scala 39:67 PEArray.scala 101:22]
  wire [2:0] _GEN_348 = _T_41 ? _GEN_331 : state; // @[Conditional.scala 39:67 PEArray.scala 100:22]
  wire [5:0] _GEN_353 = _T_31 ? _GEN_334 : _GEN_346; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_354 = _T_31 ? _GEN_330 : _GEN_347; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_355 = _T_31 ? _GEN_331 : _GEN_348; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_356 = _T_22 ? _GEN_330 : _GEN_354; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_357 = _T_22 ? _GEN_329 : _GEN_353; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_458 = _T_22 ? _GEN_331 : _GEN_355; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_690 = _T_3 ? _GEN_118 : {{2'd0}, GRU_out_width}; // @[Conditional.scala 40:58 PEArray.scala 104:26]
  FP16MulAdder FP16MAC ( // @[PEArray.scala 72:23]
    .io_a(FP16MAC_io_a),
    .io_b(FP16MAC_io_b),
    .io_c(FP16MAC_io_c),
    .io_out(FP16MAC_io_out)
  );
  assign io_ToRightPE = mux3out_reg; // @[PEArray.scala 95:16]
  assign io_ToBelowPE = mux2out_reg; // @[PEArray.scala 94:16]
  assign FP16MAC_io_a = sel1 ? io_FromL1 : io_FromLeftPE; // @[PEArray.scala 50:14 PEArray.scala 50:23 PEArray.scala 51:24]
  assign FP16MAC_io_b = sel5 ? mux4out : _GEN_105; // @[PEArray.scala 77:13 PEArray.scala 78:18 PEArray.scala 81:18]
  assign FP16MAC_io_c = sel5 ? _GEN_105 : mux4out; // @[PEArray.scala 77:13 PEArray.scala 79:18 PEArray.scala 82:18]
  always @(posedge clock) begin
    if (reset) begin // @[PEArray.scala 39:24]
      L0Index <= 6'h0; // @[PEArray.scala 39:24]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h0; // @[PEArray.scala 159:15]
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        L0Index <= 6'hc; // @[PEArray.scala 181:15]
      end else begin
        L0Index <= _GEN_357;
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_0 <= _GEN_229;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_1 <= _GEN_230;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_2 <= _GEN_231;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_3 <= _GEN_232;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_4 <= _GEN_233;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_5 <= _GEN_234;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_6 <= _GEN_235;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_7 <= _GEN_236;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_8 <= _GEN_237;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_9 <= _GEN_238;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_10 <= _GEN_239;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_11 <= _GEN_240;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_12 <= _GEN_241;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_13 <= _GEN_242;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_14 <= _GEN_243;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_15 <= _GEN_244;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_16 <= _GEN_245;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_17 <= _GEN_246;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_18 <= _GEN_247;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_19 <= _GEN_248;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_20 <= _GEN_249;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_21 <= _GEN_250;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_22 <= _GEN_251;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_23 <= _GEN_252;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_24 <= _GEN_253;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_25 <= _GEN_254;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_26 <= _GEN_255;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_27 <= _GEN_256;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_28 <= _GEN_257;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_29 <= _GEN_258;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_30 <= _GEN_259;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_31 <= _GEN_260;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_32 <= _GEN_261;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_33 <= _GEN_262;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_34 <= _GEN_263;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_35 <= _GEN_264;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_36 <= _GEN_265;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_37 <= _GEN_266;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_38 <= _GEN_267;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_39 <= _GEN_268;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_40 <= _GEN_269;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_41 <= _GEN_270;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_42 <= _GEN_271;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_43 <= _GEN_272;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_44 <= _GEN_273;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_45 <= _GEN_274;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_46 <= _GEN_275;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_47 <= _GEN_276;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_48 <= _GEN_277;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_49 <= _GEN_278;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_50 <= _GEN_279;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_51 <= _GEN_280;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_52 <= _GEN_281;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_53 <= _GEN_282;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_54 <= _GEN_283;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_55 <= _GEN_284;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_56 <= _GEN_285;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_57 <= _GEN_286;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_58 <= _GEN_287;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_59 <= _GEN_288;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_60 <= _GEN_289;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_61 <= _GEN_290;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_62 <= _GEN_291;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_63 <= _GEN_292;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_64 <= _GEN_293;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_65 <= _GEN_294;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_66 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_67 <= _GEN_296;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_68 <= _GEN_297;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_69 <= _GEN_298;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_70 <= _GEN_299;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_71 <= _GEN_300;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_72 <= _GEN_301;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_73 <= _GEN_302;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_74 <= _GEN_303;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_75 <= _GEN_304;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_76 <= _GEN_305;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_77 <= _GEN_306;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_78 <= _GEN_307;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_79 <= _GEN_308;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_80 <= _GEN_309;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_81 <= _GEN_310;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_82 <= _GEN_311;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_83 <= _GEN_312;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_84 <= _GEN_313;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_85 <= _GEN_314;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_86 <= _GEN_315;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_87 <= _GEN_316;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_88 <= _GEN_317;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_89 <= _GEN_318;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_90 <= _GEN_319;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_91 <= _GEN_320;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_92 <= _GEN_321;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_93 <= _GEN_322;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_94 <= _GEN_323;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_95 <= _GEN_324;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_96 <= _GEN_325;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_97 <= _GEN_326;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_98 <= _GEN_327;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_99 <= _GEN_328;
          end
        end
      end
    end
    if (reset) begin // @[PEArray.scala 100:22]
      state <= 3'h0; // @[PEArray.scala 100:22]
    end else if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[2]) begin // @[PEArray.scala 116:57]
        state <= 3'h1;
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      if (count == 10'h33) begin // @[PEArray.scala 164:27]
        state <= 3'h0; // @[PEArray.scala 166:15]
      end
    end else if (_T_16) begin // @[Conditional.scala 39:67]
      state <= _GEN_126;
    end else begin
      state <= _GEN_458;
    end
    if (reset) begin // @[PEArray.scala 90:28]
      mux2out_reg <= 16'h0; // @[PEArray.scala 90:28]
    end else begin
      mux2out_reg <= MAC_out; // @[PEArray.scala 90:28]
    end
    if (reset) begin // @[PEArray.scala 91:28]
      mux3out_reg <= 16'h0; // @[PEArray.scala 91:28]
    end else if (sel3) begin // @[PEArray.scala 56:14]
      mux3out_reg <= MAC_out; // @[PEArray.scala 56:23]
    end else if (sel1) begin // @[PEArray.scala 50:14]
      mux3out_reg <= io_FromL1; // @[PEArray.scala 50:23]
    end else begin
      mux3out_reg <= io_FromLeftPE; // @[PEArray.scala 51:24]
    end
    if (reset) begin // @[PEArray.scala 101:22]
      count <= 10'h0; // @[PEArray.scala 101:22]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        if (count == 10'h33) begin // @[PEArray.scala 164:27]
          count <= 10'h0; // @[PEArray.scala 165:15]
        end else begin
          count <= _GEN_120;
        end
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        count <= _GEN_125;
      end else begin
        count <= _GEN_356;
      end
    end
    GRU_out_width <= _GEN_690[5:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  L0Index = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  L0Memory_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  L0Memory_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  L0Memory_2 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  L0Memory_3 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  L0Memory_4 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  L0Memory_5 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  L0Memory_6 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  L0Memory_7 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  L0Memory_8 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  L0Memory_9 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  L0Memory_10 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  L0Memory_11 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  L0Memory_12 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  L0Memory_13 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  L0Memory_14 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  L0Memory_15 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  L0Memory_16 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  L0Memory_17 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  L0Memory_18 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  L0Memory_19 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  L0Memory_20 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  L0Memory_21 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  L0Memory_22 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  L0Memory_23 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  L0Memory_24 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  L0Memory_25 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  L0Memory_26 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  L0Memory_27 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  L0Memory_28 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  L0Memory_29 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  L0Memory_30 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  L0Memory_31 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  L0Memory_32 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  L0Memory_33 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  L0Memory_34 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  L0Memory_35 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  L0Memory_36 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  L0Memory_37 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  L0Memory_38 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  L0Memory_39 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  L0Memory_40 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  L0Memory_41 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  L0Memory_42 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  L0Memory_43 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  L0Memory_44 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  L0Memory_45 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  L0Memory_46 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  L0Memory_47 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  L0Memory_48 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  L0Memory_49 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  L0Memory_50 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  L0Memory_51 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  L0Memory_52 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  L0Memory_53 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  L0Memory_54 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  L0Memory_55 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  L0Memory_56 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  L0Memory_57 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  L0Memory_58 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  L0Memory_59 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  L0Memory_60 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  L0Memory_61 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  L0Memory_62 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  L0Memory_63 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  L0Memory_64 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  L0Memory_65 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  L0Memory_66 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  L0Memory_67 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  L0Memory_68 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  L0Memory_69 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  L0Memory_70 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  L0Memory_71 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  L0Memory_72 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  L0Memory_73 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  L0Memory_74 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  L0Memory_75 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  L0Memory_76 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  L0Memory_77 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  L0Memory_78 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  L0Memory_79 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  L0Memory_80 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  L0Memory_81 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  L0Memory_82 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  L0Memory_83 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  L0Memory_84 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  L0Memory_85 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  L0Memory_86 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  L0Memory_87 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  L0Memory_88 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  L0Memory_89 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  L0Memory_90 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  L0Memory_91 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  L0Memory_92 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  L0Memory_93 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  L0Memory_94 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  L0Memory_95 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  L0Memory_96 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  L0Memory_97 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  L0Memory_98 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  L0Memory_99 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  state = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  mux2out_reg = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  mux3out_reg = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  count = _RAND_104[9:0];
  _RAND_105 = {1{`RANDOM}};
  GRU_out_width = _RAND_105[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PE_28(
  input         clock,
  input         reset,
  input  [15:0] io_FromAbovePE,
  input  [15:0] io_FromLeftPE,
  input  [15:0] io_FromL1,
  input  [11:0] io_control_signal_mask,
  output [15:0] io_ToRightPE,
  output [15:0] io_ToBelowPE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] FP16MAC_io_a; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_b; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_c; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_out; // @[PEArray.scala 72:23]
  reg [5:0] L0Index; // @[PEArray.scala 39:24]
  reg [15:0] L0Memory_0; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_1; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_2; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_3; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_4; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_5; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_6; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_7; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_8; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_9; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_10; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_11; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_12; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_13; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_14; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_15; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_16; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_17; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_18; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_19; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_20; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_21; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_22; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_23; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_24; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_25; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_26; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_27; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_28; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_29; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_30; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_31; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_32; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_33; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_34; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_35; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_36; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_37; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_38; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_39; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_40; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_41; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_42; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_43; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_44; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_45; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_46; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_47; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_48; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_49; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_50; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_51; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_52; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_53; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_54; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_55; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_56; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_57; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_58; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_59; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_60; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_61; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_62; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_63; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_64; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_65; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_66; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_67; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_68; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_69; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_70; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_71; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_72; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_73; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_74; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_75; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_76; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_77; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_78; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_79; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_80; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_81; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_82; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_83; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_84; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_85; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_86; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_87; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_88; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_89; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_90; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_91; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_92; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_93; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_94; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_95; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_96; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_97; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_98; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_99; // @[PEArray.scala 40:21]
  reg [2:0] state; // @[PEArray.scala 100:22]
  wire  _T_3 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_12 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_16 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_22 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_31 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_41 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_342 = _T_41 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 231:12 PEArray.scala 32:8]
  wire  _GEN_349 = _T_31 ? 1'h0 : _GEN_342; // @[Conditional.scala 39:67 PEArray.scala 208:12]
  wire  _GEN_459 = _T_22 | _GEN_349; // @[Conditional.scala 39:67 PEArray.scala 32:8]
  wire  _GEN_463 = _T_16 ? 1'h0 : _GEN_459; // @[Conditional.scala 39:67]
  wire  _GEN_572 = _T_12 | _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 149:12]
  wire  sel1 = _T_3 | _GEN_572; // @[Conditional.scala 40:58 PEArray.scala 108:12]
  wire [15:0] MAC_out = FP16MAC_io_out; // @[PEArray.scala 47:21 PEArray.scala 85:11]
  wire  _GEN_465 = _T_16 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 177:12]
  wire  _GEN_580 = _T_12 | _GEN_465; // @[Conditional.scala 39:67 PEArray.scala 34:8]
  wire  sel3 = _T_3 | _GEN_580; // @[Conditional.scala 40:58 PEArray.scala 110:12]
  wire [1:0] _GEN_344 = _T_41 ? 2'h2 : 2'h0; // @[Conditional.scala 39:67 PEArray.scala 233:12 PEArray.scala 35:8]
  wire [1:0] _GEN_351 = _T_31 ? 2'h2 : _GEN_344; // @[Conditional.scala 39:67 PEArray.scala 210:12]
  wire [1:0] _GEN_461 = _T_22 ? 2'h0 : _GEN_351; // @[Conditional.scala 39:67 PEArray.scala 35:8]
  wire [1:0] _GEN_466 = _T_16 ? 2'h0 : _GEN_461; // @[Conditional.scala 39:67 PEArray.scala 178:12]
  wire [1:0] _GEN_574 = _T_12 ? 2'h1 : _GEN_466; // @[Conditional.scala 39:67]
  wire [1:0] sel4 = _T_3 ? 2'h0 : _GEN_574; // @[Conditional.scala 40:58 PEArray.scala 111:12]
  wire [15:0] _GEN_3 = sel4 == 2'h2 ? io_FromL1 : 16'h0; // @[PEArray.scala 65:28 PEArray.scala 66:15 PEArray.scala 69:15]
  wire [15:0] _GEN_4 = sel4 == 2'h1 ? io_FromAbovePE : _GEN_3; // @[PEArray.scala 62:28 PEArray.scala 63:15]
  wire [15:0] mux4out = sel4 == 2'h0 ? 16'h0 : _GEN_4; // @[PEArray.scala 59:22 PEArray.scala 60:13]
  wire [15:0] _GEN_7 = 6'h1 == L0Index ? L0Memory_1 : L0Memory_0; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_8 = 6'h2 == L0Index ? L0Memory_2 : _GEN_7; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_9 = 6'h3 == L0Index ? L0Memory_3 : _GEN_8; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_10 = 6'h4 == L0Index ? L0Memory_4 : _GEN_9; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_11 = 6'h5 == L0Index ? L0Memory_5 : _GEN_10; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_12 = 6'h6 == L0Index ? L0Memory_6 : _GEN_11; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_13 = 6'h7 == L0Index ? L0Memory_7 : _GEN_12; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_14 = 6'h8 == L0Index ? L0Memory_8 : _GEN_13; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_15 = 6'h9 == L0Index ? L0Memory_9 : _GEN_14; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_16 = 6'ha == L0Index ? L0Memory_10 : _GEN_15; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_17 = 6'hb == L0Index ? L0Memory_11 : _GEN_16; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_18 = 6'hc == L0Index ? L0Memory_12 : _GEN_17; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_19 = 6'hd == L0Index ? L0Memory_13 : _GEN_18; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_20 = 6'he == L0Index ? L0Memory_14 : _GEN_19; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_21 = 6'hf == L0Index ? L0Memory_15 : _GEN_20; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_22 = 6'h10 == L0Index ? L0Memory_16 : _GEN_21; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_23 = 6'h11 == L0Index ? L0Memory_17 : _GEN_22; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_24 = 6'h12 == L0Index ? L0Memory_18 : _GEN_23; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_25 = 6'h13 == L0Index ? L0Memory_19 : _GEN_24; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_26 = 6'h14 == L0Index ? L0Memory_20 : _GEN_25; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_27 = 6'h15 == L0Index ? L0Memory_21 : _GEN_26; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_28 = 6'h16 == L0Index ? L0Memory_22 : _GEN_27; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_29 = 6'h17 == L0Index ? L0Memory_23 : _GEN_28; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_30 = 6'h18 == L0Index ? L0Memory_24 : _GEN_29; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_31 = 6'h19 == L0Index ? L0Memory_25 : _GEN_30; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_32 = 6'h1a == L0Index ? L0Memory_26 : _GEN_31; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_33 = 6'h1b == L0Index ? L0Memory_27 : _GEN_32; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_34 = 6'h1c == L0Index ? L0Memory_28 : _GEN_33; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_35 = 6'h1d == L0Index ? L0Memory_29 : _GEN_34; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_36 = 6'h1e == L0Index ? L0Memory_30 : _GEN_35; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_37 = 6'h1f == L0Index ? L0Memory_31 : _GEN_36; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_38 = 6'h20 == L0Index ? L0Memory_32 : _GEN_37; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_39 = 6'h21 == L0Index ? L0Memory_33 : _GEN_38; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_40 = 6'h22 == L0Index ? L0Memory_34 : _GEN_39; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_41 = 6'h23 == L0Index ? L0Memory_35 : _GEN_40; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_42 = 6'h24 == L0Index ? L0Memory_36 : _GEN_41; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_43 = 6'h25 == L0Index ? L0Memory_37 : _GEN_42; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_44 = 6'h26 == L0Index ? L0Memory_38 : _GEN_43; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_45 = 6'h27 == L0Index ? L0Memory_39 : _GEN_44; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_46 = 6'h28 == L0Index ? L0Memory_40 : _GEN_45; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_47 = 6'h29 == L0Index ? L0Memory_41 : _GEN_46; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_48 = 6'h2a == L0Index ? L0Memory_42 : _GEN_47; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_49 = 6'h2b == L0Index ? L0Memory_43 : _GEN_48; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_50 = 6'h2c == L0Index ? L0Memory_44 : _GEN_49; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_51 = 6'h2d == L0Index ? L0Memory_45 : _GEN_50; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_52 = 6'h2e == L0Index ? L0Memory_46 : _GEN_51; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_53 = 6'h2f == L0Index ? L0Memory_47 : _GEN_52; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_54 = 6'h30 == L0Index ? L0Memory_48 : _GEN_53; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_55 = 6'h31 == L0Index ? L0Memory_49 : _GEN_54; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_56 = 6'h32 == L0Index ? L0Memory_50 : _GEN_55; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_57 = 6'h33 == L0Index ? L0Memory_51 : _GEN_56; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_58 = 6'h34 == L0Index ? L0Memory_52 : _GEN_57; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_59 = 6'h35 == L0Index ? L0Memory_53 : _GEN_58; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_60 = 6'h36 == L0Index ? L0Memory_54 : _GEN_59; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_61 = 6'h37 == L0Index ? L0Memory_55 : _GEN_60; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_62 = 6'h38 == L0Index ? L0Memory_56 : _GEN_61; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_63 = 6'h39 == L0Index ? L0Memory_57 : _GEN_62; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_64 = 6'h3a == L0Index ? L0Memory_58 : _GEN_63; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_65 = 6'h3b == L0Index ? L0Memory_59 : _GEN_64; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_66 = 6'h3c == L0Index ? L0Memory_60 : _GEN_65; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_67 = 6'h3d == L0Index ? L0Memory_61 : _GEN_66; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_68 = 6'h3e == L0Index ? L0Memory_62 : _GEN_67; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_69 = 6'h3f == L0Index ? L0Memory_63 : _GEN_68; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [6:0] _GEN_793 = {{1'd0}, L0Index}; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_70 = 7'h40 == _GEN_793 ? L0Memory_64 : _GEN_69; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_71 = 7'h41 == _GEN_793 ? L0Memory_65 : _GEN_70; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_72 = 7'h42 == _GEN_793 ? L0Memory_66 : _GEN_71; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_73 = 7'h43 == _GEN_793 ? L0Memory_67 : _GEN_72; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_74 = 7'h44 == _GEN_793 ? L0Memory_68 : _GEN_73; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_75 = 7'h45 == _GEN_793 ? L0Memory_69 : _GEN_74; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_76 = 7'h46 == _GEN_793 ? L0Memory_70 : _GEN_75; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_77 = 7'h47 == _GEN_793 ? L0Memory_71 : _GEN_76; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_78 = 7'h48 == _GEN_793 ? L0Memory_72 : _GEN_77; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_79 = 7'h49 == _GEN_793 ? L0Memory_73 : _GEN_78; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_80 = 7'h4a == _GEN_793 ? L0Memory_74 : _GEN_79; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_81 = 7'h4b == _GEN_793 ? L0Memory_75 : _GEN_80; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_82 = 7'h4c == _GEN_793 ? L0Memory_76 : _GEN_81; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_83 = 7'h4d == _GEN_793 ? L0Memory_77 : _GEN_82; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_84 = 7'h4e == _GEN_793 ? L0Memory_78 : _GEN_83; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_85 = 7'h4f == _GEN_793 ? L0Memory_79 : _GEN_84; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_86 = 7'h50 == _GEN_793 ? L0Memory_80 : _GEN_85; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_87 = 7'h51 == _GEN_793 ? L0Memory_81 : _GEN_86; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_88 = 7'h52 == _GEN_793 ? L0Memory_82 : _GEN_87; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_89 = 7'h53 == _GEN_793 ? L0Memory_83 : _GEN_88; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_90 = 7'h54 == _GEN_793 ? L0Memory_84 : _GEN_89; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_91 = 7'h55 == _GEN_793 ? L0Memory_85 : _GEN_90; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_92 = 7'h56 == _GEN_793 ? L0Memory_86 : _GEN_91; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_93 = 7'h57 == _GEN_793 ? L0Memory_87 : _GEN_92; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_94 = 7'h58 == _GEN_793 ? L0Memory_88 : _GEN_93; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_95 = 7'h59 == _GEN_793 ? L0Memory_89 : _GEN_94; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_96 = 7'h5a == _GEN_793 ? L0Memory_90 : _GEN_95; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_97 = 7'h5b == _GEN_793 ? L0Memory_91 : _GEN_96; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_98 = 7'h5c == _GEN_793 ? L0Memory_92 : _GEN_97; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_99 = 7'h5d == _GEN_793 ? L0Memory_93 : _GEN_98; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_100 = 7'h5e == _GEN_793 ? L0Memory_94 : _GEN_99; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_101 = 7'h5f == _GEN_793 ? L0Memory_95 : _GEN_100; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_102 = 7'h60 == _GEN_793 ? L0Memory_96 : _GEN_101; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_103 = 7'h61 == _GEN_793 ? L0Memory_97 : _GEN_102; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_104 = 7'h62 == _GEN_793 ? L0Memory_98 : _GEN_103; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_105 = 7'h63 == _GEN_793 ? L0Memory_99 : _GEN_104; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire  _GEN_575 = _T_12 ? 1'h0 : _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 157:12]
  wire  sel5 = _T_3 ? 1'h0 : _GEN_575; // @[Conditional.scala 40:58 PEArray.scala 112:12]
  reg [15:0] mux2out_reg; // @[PEArray.scala 90:28]
  reg [15:0] mux3out_reg; // @[PEArray.scala 91:28]
  reg [9:0] count; // @[PEArray.scala 101:22]
  reg [5:0] GRU_out_width; // @[PEArray.scala 104:26]
  wire [7:0] _GEN_118 = io_control_signal_mask[2] ? 8'h0 : {{2'd0}, GRU_out_width}; // @[PEArray.scala 116:57 PEArray.scala 145:23 PEArray.scala 104:26]
  wire [9:0] _count_T_1 = count + 10'h1; // @[PEArray.scala 162:24]
  wire [9:0] _GEN_120 = count != 10'h33 ? _count_T_1 : count; // @[PEArray.scala 161:27 PEArray.scala 162:15 PEArray.scala 101:22]
  wire [9:0] _GEN_124 = count != 10'h188 ? _count_T_1 : count; // @[PEArray.scala 183:28 PEArray.scala 184:15 PEArray.scala 101:22]
  wire [9:0] _GEN_125 = count == 10'h188 ? 10'h0 : _GEN_124; // @[PEArray.scala 186:28 PEArray.scala 187:15]
  wire [2:0] _GEN_126 = count == 10'h188 ? 3'h0 : state; // @[PEArray.scala 186:28 PEArray.scala 188:15 PEArray.scala 100:22]
  wire [9:0] _GEN_127 = count != 10'h0 ? _count_T_1 : count; // @[PEArray.scala 192:32 PEArray.scala 193:15 PEArray.scala 101:22]
  wire  _T_24 = count == 10'h0; // @[PEArray.scala 195:18]
  wire [5:0] _GEN_128 = count == 10'h0 ? 6'h0 : L0Index; // @[PEArray.scala 195:26 PEArray.scala 196:17 PEArray.scala 39:24]
  wire [9:0] _T_27 = 10'h0 - 10'h1; // @[PEArray.scala 198:51]
  wire [15:0] _GEN_129 = 6'h0 == L0Index ? io_FromL1 : L0Memory_0; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_130 = 6'h1 == L0Index ? io_FromL1 : L0Memory_1; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_131 = 6'h2 == L0Index ? io_FromL1 : L0Memory_2; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_132 = 6'h3 == L0Index ? io_FromL1 : L0Memory_3; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_133 = 6'h4 == L0Index ? io_FromL1 : L0Memory_4; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_134 = 6'h5 == L0Index ? io_FromL1 : L0Memory_5; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_135 = 6'h6 == L0Index ? io_FromL1 : L0Memory_6; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_136 = 6'h7 == L0Index ? io_FromL1 : L0Memory_7; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_137 = 6'h8 == L0Index ? io_FromL1 : L0Memory_8; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_138 = 6'h9 == L0Index ? io_FromL1 : L0Memory_9; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_139 = 6'ha == L0Index ? io_FromL1 : L0Memory_10; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_140 = 6'hb == L0Index ? io_FromL1 : L0Memory_11; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_141 = 6'hc == L0Index ? io_FromL1 : L0Memory_12; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_142 = 6'hd == L0Index ? io_FromL1 : L0Memory_13; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_143 = 6'he == L0Index ? io_FromL1 : L0Memory_14; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_144 = 6'hf == L0Index ? io_FromL1 : L0Memory_15; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_145 = 6'h10 == L0Index ? io_FromL1 : L0Memory_16; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_146 = 6'h11 == L0Index ? io_FromL1 : L0Memory_17; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_147 = 6'h12 == L0Index ? io_FromL1 : L0Memory_18; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_148 = 6'h13 == L0Index ? io_FromL1 : L0Memory_19; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_149 = 6'h14 == L0Index ? io_FromL1 : L0Memory_20; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_150 = 6'h15 == L0Index ? io_FromL1 : L0Memory_21; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_151 = 6'h16 == L0Index ? io_FromL1 : L0Memory_22; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_152 = 6'h17 == L0Index ? io_FromL1 : L0Memory_23; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_153 = 6'h18 == L0Index ? io_FromL1 : L0Memory_24; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_154 = 6'h19 == L0Index ? io_FromL1 : L0Memory_25; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_155 = 6'h1a == L0Index ? io_FromL1 : L0Memory_26; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_156 = 6'h1b == L0Index ? io_FromL1 : L0Memory_27; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_157 = 6'h1c == L0Index ? io_FromL1 : L0Memory_28; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_158 = 6'h1d == L0Index ? io_FromL1 : L0Memory_29; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_159 = 6'h1e == L0Index ? io_FromL1 : L0Memory_30; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_160 = 6'h1f == L0Index ? io_FromL1 : L0Memory_31; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_161 = 6'h20 == L0Index ? io_FromL1 : L0Memory_32; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_162 = 6'h21 == L0Index ? io_FromL1 : L0Memory_33; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_163 = 6'h22 == L0Index ? io_FromL1 : L0Memory_34; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_164 = 6'h23 == L0Index ? io_FromL1 : L0Memory_35; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_165 = 6'h24 == L0Index ? io_FromL1 : L0Memory_36; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_166 = 6'h25 == L0Index ? io_FromL1 : L0Memory_37; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_167 = 6'h26 == L0Index ? io_FromL1 : L0Memory_38; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_168 = 6'h27 == L0Index ? io_FromL1 : L0Memory_39; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_169 = 6'h28 == L0Index ? io_FromL1 : L0Memory_40; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_170 = 6'h29 == L0Index ? io_FromL1 : L0Memory_41; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_171 = 6'h2a == L0Index ? io_FromL1 : L0Memory_42; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_172 = 6'h2b == L0Index ? io_FromL1 : L0Memory_43; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_173 = 6'h2c == L0Index ? io_FromL1 : L0Memory_44; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_174 = 6'h2d == L0Index ? io_FromL1 : L0Memory_45; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_175 = 6'h2e == L0Index ? io_FromL1 : L0Memory_46; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_176 = 6'h2f == L0Index ? io_FromL1 : L0Memory_47; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_177 = 6'h30 == L0Index ? io_FromL1 : L0Memory_48; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_178 = 6'h31 == L0Index ? io_FromL1 : L0Memory_49; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_179 = 6'h32 == L0Index ? io_FromL1 : L0Memory_50; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_180 = 6'h33 == L0Index ? io_FromL1 : L0Memory_51; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_181 = 6'h34 == L0Index ? io_FromL1 : L0Memory_52; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_182 = 6'h35 == L0Index ? io_FromL1 : L0Memory_53; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_183 = 6'h36 == L0Index ? io_FromL1 : L0Memory_54; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_184 = 6'h37 == L0Index ? io_FromL1 : L0Memory_55; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_185 = 6'h38 == L0Index ? io_FromL1 : L0Memory_56; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_186 = 6'h39 == L0Index ? io_FromL1 : L0Memory_57; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_187 = 6'h3a == L0Index ? io_FromL1 : L0Memory_58; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_188 = 6'h3b == L0Index ? io_FromL1 : L0Memory_59; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_189 = 6'h3c == L0Index ? io_FromL1 : L0Memory_60; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_190 = 6'h3d == L0Index ? io_FromL1 : L0Memory_61; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_191 = 6'h3e == L0Index ? io_FromL1 : L0Memory_62; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_192 = 6'h3f == L0Index ? io_FromL1 : L0Memory_63; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_193 = 7'h40 == _GEN_793 ? io_FromL1 : L0Memory_64; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_194 = 7'h41 == _GEN_793 ? io_FromL1 : L0Memory_65; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_195 = 7'h42 == _GEN_793 ? io_FromL1 : L0Memory_66; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_196 = 7'h43 == _GEN_793 ? io_FromL1 : L0Memory_67; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_197 = 7'h44 == _GEN_793 ? io_FromL1 : L0Memory_68; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_198 = 7'h45 == _GEN_793 ? io_FromL1 : L0Memory_69; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_199 = 7'h46 == _GEN_793 ? io_FromL1 : L0Memory_70; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_200 = 7'h47 == _GEN_793 ? io_FromL1 : L0Memory_71; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_201 = 7'h48 == _GEN_793 ? io_FromL1 : L0Memory_72; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_202 = 7'h49 == _GEN_793 ? io_FromL1 : L0Memory_73; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_203 = 7'h4a == _GEN_793 ? io_FromL1 : L0Memory_74; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_204 = 7'h4b == _GEN_793 ? io_FromL1 : L0Memory_75; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_205 = 7'h4c == _GEN_793 ? io_FromL1 : L0Memory_76; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_206 = 7'h4d == _GEN_793 ? io_FromL1 : L0Memory_77; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_207 = 7'h4e == _GEN_793 ? io_FromL1 : L0Memory_78; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_208 = 7'h4f == _GEN_793 ? io_FromL1 : L0Memory_79; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_209 = 7'h50 == _GEN_793 ? io_FromL1 : L0Memory_80; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_210 = 7'h51 == _GEN_793 ? io_FromL1 : L0Memory_81; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_211 = 7'h52 == _GEN_793 ? io_FromL1 : L0Memory_82; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_212 = 7'h53 == _GEN_793 ? io_FromL1 : L0Memory_83; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_213 = 7'h54 == _GEN_793 ? io_FromL1 : L0Memory_84; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_214 = 7'h55 == _GEN_793 ? io_FromL1 : L0Memory_85; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_215 = 7'h56 == _GEN_793 ? io_FromL1 : L0Memory_86; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_216 = 7'h57 == _GEN_793 ? io_FromL1 : L0Memory_87; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_217 = 7'h58 == _GEN_793 ? io_FromL1 : L0Memory_88; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_218 = 7'h59 == _GEN_793 ? io_FromL1 : L0Memory_89; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_219 = 7'h5a == _GEN_793 ? io_FromL1 : L0Memory_90; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_220 = 7'h5b == _GEN_793 ? io_FromL1 : L0Memory_91; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_221 = 7'h5c == _GEN_793 ? io_FromL1 : L0Memory_92; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_222 = 7'h5d == _GEN_793 ? io_FromL1 : L0Memory_93; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_223 = 7'h5e == _GEN_793 ? io_FromL1 : L0Memory_94; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_224 = 7'h5f == _GEN_793 ? io_FromL1 : L0Memory_95; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_225 = 7'h60 == _GEN_793 ? io_FromL1 : L0Memory_96; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_226 = 7'h61 == _GEN_793 ? io_FromL1 : L0Memory_97; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_227 = 7'h62 == _GEN_793 ? io_FromL1 : L0Memory_98; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_228 = 7'h63 == _GEN_793 ? io_FromL1 : L0Memory_99; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [5:0] _L0Index_T_2 = L0Index + 6'h1; // @[PEArray.scala 200:28]
  wire [15:0] _GEN_229 = count >= 10'h1 & count <= _T_27 ? _GEN_129 : L0Memory_0; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_230 = count >= 10'h1 & count <= _T_27 ? _GEN_130 : L0Memory_1; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_231 = count >= 10'h1 & count <= _T_27 ? _GEN_131 : L0Memory_2; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_232 = count >= 10'h1 & count <= _T_27 ? _GEN_132 : L0Memory_3; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_233 = count >= 10'h1 & count <= _T_27 ? _GEN_133 : L0Memory_4; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_234 = count >= 10'h1 & count <= _T_27 ? _GEN_134 : L0Memory_5; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_235 = count >= 10'h1 & count <= _T_27 ? _GEN_135 : L0Memory_6; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_236 = count >= 10'h1 & count <= _T_27 ? _GEN_136 : L0Memory_7; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_237 = count >= 10'h1 & count <= _T_27 ? _GEN_137 : L0Memory_8; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_238 = count >= 10'h1 & count <= _T_27 ? _GEN_138 : L0Memory_9; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_239 = count >= 10'h1 & count <= _T_27 ? _GEN_139 : L0Memory_10; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_240 = count >= 10'h1 & count <= _T_27 ? _GEN_140 : L0Memory_11; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_241 = count >= 10'h1 & count <= _T_27 ? _GEN_141 : L0Memory_12; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_242 = count >= 10'h1 & count <= _T_27 ? _GEN_142 : L0Memory_13; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_243 = count >= 10'h1 & count <= _T_27 ? _GEN_143 : L0Memory_14; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_244 = count >= 10'h1 & count <= _T_27 ? _GEN_144 : L0Memory_15; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_245 = count >= 10'h1 & count <= _T_27 ? _GEN_145 : L0Memory_16; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_246 = count >= 10'h1 & count <= _T_27 ? _GEN_146 : L0Memory_17; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_247 = count >= 10'h1 & count <= _T_27 ? _GEN_147 : L0Memory_18; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_248 = count >= 10'h1 & count <= _T_27 ? _GEN_148 : L0Memory_19; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_249 = count >= 10'h1 & count <= _T_27 ? _GEN_149 : L0Memory_20; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_250 = count >= 10'h1 & count <= _T_27 ? _GEN_150 : L0Memory_21; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_251 = count >= 10'h1 & count <= _T_27 ? _GEN_151 : L0Memory_22; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_252 = count >= 10'h1 & count <= _T_27 ? _GEN_152 : L0Memory_23; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_253 = count >= 10'h1 & count <= _T_27 ? _GEN_153 : L0Memory_24; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_254 = count >= 10'h1 & count <= _T_27 ? _GEN_154 : L0Memory_25; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_255 = count >= 10'h1 & count <= _T_27 ? _GEN_155 : L0Memory_26; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_256 = count >= 10'h1 & count <= _T_27 ? _GEN_156 : L0Memory_27; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_257 = count >= 10'h1 & count <= _T_27 ? _GEN_157 : L0Memory_28; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_258 = count >= 10'h1 & count <= _T_27 ? _GEN_158 : L0Memory_29; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_259 = count >= 10'h1 & count <= _T_27 ? _GEN_159 : L0Memory_30; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_260 = count >= 10'h1 & count <= _T_27 ? _GEN_160 : L0Memory_31; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_261 = count >= 10'h1 & count <= _T_27 ? _GEN_161 : L0Memory_32; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_262 = count >= 10'h1 & count <= _T_27 ? _GEN_162 : L0Memory_33; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_263 = count >= 10'h1 & count <= _T_27 ? _GEN_163 : L0Memory_34; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_264 = count >= 10'h1 & count <= _T_27 ? _GEN_164 : L0Memory_35; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_265 = count >= 10'h1 & count <= _T_27 ? _GEN_165 : L0Memory_36; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_266 = count >= 10'h1 & count <= _T_27 ? _GEN_166 : L0Memory_37; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_267 = count >= 10'h1 & count <= _T_27 ? _GEN_167 : L0Memory_38; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_268 = count >= 10'h1 & count <= _T_27 ? _GEN_168 : L0Memory_39; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_269 = count >= 10'h1 & count <= _T_27 ? _GEN_169 : L0Memory_40; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_270 = count >= 10'h1 & count <= _T_27 ? _GEN_170 : L0Memory_41; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_271 = count >= 10'h1 & count <= _T_27 ? _GEN_171 : L0Memory_42; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_272 = count >= 10'h1 & count <= _T_27 ? _GEN_172 : L0Memory_43; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_273 = count >= 10'h1 & count <= _T_27 ? _GEN_173 : L0Memory_44; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_274 = count >= 10'h1 & count <= _T_27 ? _GEN_174 : L0Memory_45; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_275 = count >= 10'h1 & count <= _T_27 ? _GEN_175 : L0Memory_46; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_276 = count >= 10'h1 & count <= _T_27 ? _GEN_176 : L0Memory_47; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_277 = count >= 10'h1 & count <= _T_27 ? _GEN_177 : L0Memory_48; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_278 = count >= 10'h1 & count <= _T_27 ? _GEN_178 : L0Memory_49; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_279 = count >= 10'h1 & count <= _T_27 ? _GEN_179 : L0Memory_50; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_280 = count >= 10'h1 & count <= _T_27 ? _GEN_180 : L0Memory_51; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_281 = count >= 10'h1 & count <= _T_27 ? _GEN_181 : L0Memory_52; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_282 = count >= 10'h1 & count <= _T_27 ? _GEN_182 : L0Memory_53; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_283 = count >= 10'h1 & count <= _T_27 ? _GEN_183 : L0Memory_54; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_284 = count >= 10'h1 & count <= _T_27 ? _GEN_184 : L0Memory_55; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_285 = count >= 10'h1 & count <= _T_27 ? _GEN_185 : L0Memory_56; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_286 = count >= 10'h1 & count <= _T_27 ? _GEN_186 : L0Memory_57; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_287 = count >= 10'h1 & count <= _T_27 ? _GEN_187 : L0Memory_58; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_288 = count >= 10'h1 & count <= _T_27 ? _GEN_188 : L0Memory_59; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_289 = count >= 10'h1 & count <= _T_27 ? _GEN_189 : L0Memory_60; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_290 = count >= 10'h1 & count <= _T_27 ? _GEN_190 : L0Memory_61; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_291 = count >= 10'h1 & count <= _T_27 ? _GEN_191 : L0Memory_62; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_292 = count >= 10'h1 & count <= _T_27 ? _GEN_192 : L0Memory_63; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_293 = count >= 10'h1 & count <= _T_27 ? _GEN_193 : L0Memory_64; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_294 = count >= 10'h1 & count <= _T_27 ? _GEN_194 : L0Memory_65; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_295 = count >= 10'h1 & count <= _T_27 ? _GEN_195 : L0Memory_66; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_296 = count >= 10'h1 & count <= _T_27 ? _GEN_196 : L0Memory_67; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_297 = count >= 10'h1 & count <= _T_27 ? _GEN_197 : L0Memory_68; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_298 = count >= 10'h1 & count <= _T_27 ? _GEN_198 : L0Memory_69; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_299 = count >= 10'h1 & count <= _T_27 ? _GEN_199 : L0Memory_70; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_300 = count >= 10'h1 & count <= _T_27 ? _GEN_200 : L0Memory_71; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_301 = count >= 10'h1 & count <= _T_27 ? _GEN_201 : L0Memory_72; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_302 = count >= 10'h1 & count <= _T_27 ? _GEN_202 : L0Memory_73; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_303 = count >= 10'h1 & count <= _T_27 ? _GEN_203 : L0Memory_74; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_304 = count >= 10'h1 & count <= _T_27 ? _GEN_204 : L0Memory_75; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_305 = count >= 10'h1 & count <= _T_27 ? _GEN_205 : L0Memory_76; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_306 = count >= 10'h1 & count <= _T_27 ? _GEN_206 : L0Memory_77; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_307 = count >= 10'h1 & count <= _T_27 ? _GEN_207 : L0Memory_78; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_308 = count >= 10'h1 & count <= _T_27 ? _GEN_208 : L0Memory_79; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_309 = count >= 10'h1 & count <= _T_27 ? _GEN_209 : L0Memory_80; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_310 = count >= 10'h1 & count <= _T_27 ? _GEN_210 : L0Memory_81; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_311 = count >= 10'h1 & count <= _T_27 ? _GEN_211 : L0Memory_82; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_312 = count >= 10'h1 & count <= _T_27 ? _GEN_212 : L0Memory_83; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_313 = count >= 10'h1 & count <= _T_27 ? _GEN_213 : L0Memory_84; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_314 = count >= 10'h1 & count <= _T_27 ? _GEN_214 : L0Memory_85; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_315 = count >= 10'h1 & count <= _T_27 ? _GEN_215 : L0Memory_86; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_316 = count >= 10'h1 & count <= _T_27 ? _GEN_216 : L0Memory_87; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_317 = count >= 10'h1 & count <= _T_27 ? _GEN_217 : L0Memory_88; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_318 = count >= 10'h1 & count <= _T_27 ? _GEN_218 : L0Memory_89; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_319 = count >= 10'h1 & count <= _T_27 ? _GEN_219 : L0Memory_90; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_320 = count >= 10'h1 & count <= _T_27 ? _GEN_220 : L0Memory_91; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_321 = count >= 10'h1 & count <= _T_27 ? _GEN_221 : L0Memory_92; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_322 = count >= 10'h1 & count <= _T_27 ? _GEN_222 : L0Memory_93; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_323 = count >= 10'h1 & count <= _T_27 ? _GEN_223 : L0Memory_94; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_324 = count >= 10'h1 & count <= _T_27 ? _GEN_224 : L0Memory_95; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_325 = count >= 10'h1 & count <= _T_27 ? _GEN_225 : L0Memory_96; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_326 = count >= 10'h1 & count <= _T_27 ? _GEN_226 : L0Memory_97; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_327 = count >= 10'h1 & count <= _T_27 ? _GEN_227 : L0Memory_98; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_328 = count >= 10'h1 & count <= _T_27 ? _GEN_228 : L0Memory_99; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [5:0] _GEN_329 = count >= 10'h1 & count <= _T_27 ? _L0Index_T_2 : _GEN_128; // @[PEArray.scala 198:59 PEArray.scala 200:17]
  wire [9:0] _GEN_330 = _T_24 ? 10'h0 : _GEN_127; // @[PEArray.scala 202:32 PEArray.scala 203:15]
  wire [2:0] _GEN_331 = _T_24 ? 3'h0 : state; // @[PEArray.scala 202:32 PEArray.scala 204:15 PEArray.scala 100:22]
  wire [9:0] _GEN_865 = {{4'd0}, GRU_out_width}; // @[PEArray.scala 220:19]
  wire [9:0] _GEN_0 = count % _GEN_865; // @[PEArray.scala 220:19]
  wire [5:0] _T_36 = _GEN_0[5:0]; // @[PEArray.scala 220:19]
  wire [5:0] _T_38 = GRU_out_width - 6'h1; // @[PEArray.scala 220:55]
  wire [5:0] _GEN_334 = _T_36 == _T_38 ? _L0Index_T_2 : 6'h0; // @[PEArray.scala 220:62 PEArray.scala 221:17 PEArray.scala 214:15]
  wire [5:0] _GEN_346 = _T_41 ? _GEN_334 : L0Index; // @[Conditional.scala 39:67 PEArray.scala 39:24]
  wire [9:0] _GEN_347 = _T_41 ? _GEN_330 : count; // @[Conditional.scala 39:67 PEArray.scala 101:22]
  wire [2:0] _GEN_348 = _T_41 ? _GEN_331 : state; // @[Conditional.scala 39:67 PEArray.scala 100:22]
  wire [5:0] _GEN_353 = _T_31 ? _GEN_334 : _GEN_346; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_354 = _T_31 ? _GEN_330 : _GEN_347; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_355 = _T_31 ? _GEN_331 : _GEN_348; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_356 = _T_22 ? _GEN_330 : _GEN_354; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_357 = _T_22 ? _GEN_329 : _GEN_353; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_458 = _T_22 ? _GEN_331 : _GEN_355; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_690 = _T_3 ? _GEN_118 : {{2'd0}, GRU_out_width}; // @[Conditional.scala 40:58 PEArray.scala 104:26]
  FP16MulAdder FP16MAC ( // @[PEArray.scala 72:23]
    .io_a(FP16MAC_io_a),
    .io_b(FP16MAC_io_b),
    .io_c(FP16MAC_io_c),
    .io_out(FP16MAC_io_out)
  );
  assign io_ToRightPE = mux3out_reg; // @[PEArray.scala 95:16]
  assign io_ToBelowPE = mux2out_reg; // @[PEArray.scala 94:16]
  assign FP16MAC_io_a = sel1 ? io_FromL1 : io_FromLeftPE; // @[PEArray.scala 50:14 PEArray.scala 50:23 PEArray.scala 51:24]
  assign FP16MAC_io_b = sel5 ? mux4out : _GEN_105; // @[PEArray.scala 77:13 PEArray.scala 78:18 PEArray.scala 81:18]
  assign FP16MAC_io_c = sel5 ? _GEN_105 : mux4out; // @[PEArray.scala 77:13 PEArray.scala 79:18 PEArray.scala 82:18]
  always @(posedge clock) begin
    if (reset) begin // @[PEArray.scala 39:24]
      L0Index <= 6'h0; // @[PEArray.scala 39:24]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h1; // @[PEArray.scala 159:15]
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        L0Index <= 6'hc; // @[PEArray.scala 181:15]
      end else begin
        L0Index <= _GEN_357;
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_0 <= _GEN_229;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_1 <= _GEN_230;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_2 <= _GEN_231;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_3 <= _GEN_232;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_4 <= _GEN_233;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_5 <= _GEN_234;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_6 <= _GEN_235;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_7 <= _GEN_236;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_8 <= _GEN_237;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_9 <= _GEN_238;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_10 <= _GEN_239;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_11 <= _GEN_240;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_12 <= _GEN_241;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_13 <= _GEN_242;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_14 <= _GEN_243;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_15 <= _GEN_244;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_16 <= _GEN_245;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_17 <= _GEN_246;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_18 <= _GEN_247;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_19 <= _GEN_248;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_20 <= _GEN_249;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_21 <= _GEN_250;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_22 <= _GEN_251;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_23 <= _GEN_252;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_24 <= _GEN_253;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_25 <= _GEN_254;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_26 <= _GEN_255;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_27 <= _GEN_256;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_28 <= _GEN_257;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_29 <= _GEN_258;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_30 <= _GEN_259;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_31 <= _GEN_260;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_32 <= _GEN_261;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_33 <= _GEN_262;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_34 <= _GEN_263;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_35 <= _GEN_264;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_36 <= _GEN_265;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_37 <= _GEN_266;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_38 <= _GEN_267;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_39 <= _GEN_268;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_40 <= _GEN_269;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_41 <= _GEN_270;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_42 <= _GEN_271;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_43 <= _GEN_272;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_44 <= _GEN_273;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_45 <= _GEN_274;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_46 <= _GEN_275;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_47 <= _GEN_276;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_48 <= _GEN_277;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_49 <= _GEN_278;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_50 <= _GEN_279;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_51 <= _GEN_280;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_52 <= _GEN_281;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_53 <= _GEN_282;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_54 <= _GEN_283;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_55 <= _GEN_284;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_56 <= _GEN_285;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_57 <= _GEN_286;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_58 <= _GEN_287;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_59 <= _GEN_288;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_60 <= _GEN_289;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_61 <= _GEN_290;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_62 <= _GEN_291;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_63 <= _GEN_292;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_64 <= _GEN_293;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_65 <= _GEN_294;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_66 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_67 <= _GEN_296;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_68 <= _GEN_297;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_69 <= _GEN_298;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_70 <= _GEN_299;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_71 <= _GEN_300;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_72 <= _GEN_301;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_73 <= _GEN_302;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_74 <= _GEN_303;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_75 <= _GEN_304;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_76 <= _GEN_305;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_77 <= _GEN_306;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_78 <= _GEN_307;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_79 <= _GEN_308;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_80 <= _GEN_309;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_81 <= _GEN_310;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_82 <= _GEN_311;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_83 <= _GEN_312;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_84 <= _GEN_313;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_85 <= _GEN_314;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_86 <= _GEN_315;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_87 <= _GEN_316;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_88 <= _GEN_317;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_89 <= _GEN_318;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_90 <= _GEN_319;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_91 <= _GEN_320;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_92 <= _GEN_321;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_93 <= _GEN_322;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_94 <= _GEN_323;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_95 <= _GEN_324;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_96 <= _GEN_325;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_97 <= _GEN_326;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_98 <= _GEN_327;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_99 <= _GEN_328;
          end
        end
      end
    end
    if (reset) begin // @[PEArray.scala 100:22]
      state <= 3'h0; // @[PEArray.scala 100:22]
    end else if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[2]) begin // @[PEArray.scala 116:57]
        state <= 3'h1;
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      if (count == 10'h33) begin // @[PEArray.scala 164:27]
        state <= 3'h0; // @[PEArray.scala 166:15]
      end
    end else if (_T_16) begin // @[Conditional.scala 39:67]
      state <= _GEN_126;
    end else begin
      state <= _GEN_458;
    end
    if (reset) begin // @[PEArray.scala 90:28]
      mux2out_reg <= 16'h0; // @[PEArray.scala 90:28]
    end else begin
      mux2out_reg <= MAC_out; // @[PEArray.scala 90:28]
    end
    if (reset) begin // @[PEArray.scala 91:28]
      mux3out_reg <= 16'h0; // @[PEArray.scala 91:28]
    end else if (sel3) begin // @[PEArray.scala 56:14]
      mux3out_reg <= MAC_out; // @[PEArray.scala 56:23]
    end else if (sel1) begin // @[PEArray.scala 50:14]
      mux3out_reg <= io_FromL1; // @[PEArray.scala 50:23]
    end else begin
      mux3out_reg <= io_FromLeftPE; // @[PEArray.scala 51:24]
    end
    if (reset) begin // @[PEArray.scala 101:22]
      count <= 10'h0; // @[PEArray.scala 101:22]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        if (count == 10'h33) begin // @[PEArray.scala 164:27]
          count <= 10'h0; // @[PEArray.scala 165:15]
        end else begin
          count <= _GEN_120;
        end
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        count <= _GEN_125;
      end else begin
        count <= _GEN_356;
      end
    end
    GRU_out_width <= _GEN_690[5:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  L0Index = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  L0Memory_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  L0Memory_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  L0Memory_2 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  L0Memory_3 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  L0Memory_4 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  L0Memory_5 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  L0Memory_6 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  L0Memory_7 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  L0Memory_8 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  L0Memory_9 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  L0Memory_10 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  L0Memory_11 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  L0Memory_12 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  L0Memory_13 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  L0Memory_14 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  L0Memory_15 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  L0Memory_16 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  L0Memory_17 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  L0Memory_18 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  L0Memory_19 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  L0Memory_20 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  L0Memory_21 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  L0Memory_22 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  L0Memory_23 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  L0Memory_24 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  L0Memory_25 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  L0Memory_26 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  L0Memory_27 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  L0Memory_28 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  L0Memory_29 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  L0Memory_30 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  L0Memory_31 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  L0Memory_32 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  L0Memory_33 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  L0Memory_34 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  L0Memory_35 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  L0Memory_36 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  L0Memory_37 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  L0Memory_38 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  L0Memory_39 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  L0Memory_40 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  L0Memory_41 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  L0Memory_42 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  L0Memory_43 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  L0Memory_44 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  L0Memory_45 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  L0Memory_46 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  L0Memory_47 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  L0Memory_48 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  L0Memory_49 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  L0Memory_50 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  L0Memory_51 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  L0Memory_52 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  L0Memory_53 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  L0Memory_54 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  L0Memory_55 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  L0Memory_56 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  L0Memory_57 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  L0Memory_58 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  L0Memory_59 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  L0Memory_60 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  L0Memory_61 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  L0Memory_62 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  L0Memory_63 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  L0Memory_64 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  L0Memory_65 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  L0Memory_66 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  L0Memory_67 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  L0Memory_68 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  L0Memory_69 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  L0Memory_70 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  L0Memory_71 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  L0Memory_72 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  L0Memory_73 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  L0Memory_74 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  L0Memory_75 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  L0Memory_76 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  L0Memory_77 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  L0Memory_78 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  L0Memory_79 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  L0Memory_80 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  L0Memory_81 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  L0Memory_82 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  L0Memory_83 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  L0Memory_84 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  L0Memory_85 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  L0Memory_86 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  L0Memory_87 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  L0Memory_88 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  L0Memory_89 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  L0Memory_90 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  L0Memory_91 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  L0Memory_92 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  L0Memory_93 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  L0Memory_94 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  L0Memory_95 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  L0Memory_96 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  L0Memory_97 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  L0Memory_98 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  L0Memory_99 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  state = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  mux2out_reg = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  mux3out_reg = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  count = _RAND_104[9:0];
  _RAND_105 = {1{`RANDOM}};
  GRU_out_width = _RAND_105[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PE_29(
  input         clock,
  input         reset,
  input  [15:0] io_FromAbovePE,
  input  [15:0] io_FromLeftPE,
  input  [15:0] io_FromL1,
  input  [2:0]  io_control_signal_control,
  input  [9:0]  io_control_signal_count,
  input  [5:0]  io_control_signal_L0index,
  input  [11:0] io_control_signal_mask,
  input  [7:0]  io_control_signal_gru_out_width,
  output [15:0] io_ToRightPE,
  output [15:0] io_ToBelowPE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] FP16MAC_io_a; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_b; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_c; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_out; // @[PEArray.scala 72:23]
  reg [5:0] L0Index; // @[PEArray.scala 39:24]
  reg [15:0] L0Memory_0; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_1; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_2; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_3; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_4; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_5; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_6; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_7; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_8; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_9; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_10; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_11; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_12; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_13; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_14; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_15; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_16; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_17; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_18; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_19; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_20; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_21; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_22; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_23; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_24; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_25; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_26; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_27; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_28; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_29; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_30; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_31; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_32; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_33; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_34; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_35; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_36; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_37; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_38; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_39; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_40; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_41; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_42; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_43; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_44; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_45; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_46; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_47; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_48; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_49; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_50; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_51; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_52; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_53; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_54; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_55; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_56; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_57; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_58; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_59; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_60; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_61; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_62; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_63; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_64; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_65; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_66; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_67; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_68; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_69; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_70; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_71; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_72; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_73; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_74; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_75; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_76; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_77; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_78; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_79; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_80; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_81; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_82; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_83; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_84; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_85; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_86; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_87; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_88; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_89; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_90; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_91; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_92; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_93; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_94; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_95; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_96; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_97; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_98; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_99; // @[PEArray.scala 40:21]
  reg [2:0] state; // @[PEArray.scala 100:22]
  wire  _T_3 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_12 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_16 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_22 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_31 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_41 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_342 = _T_41 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 231:12 PEArray.scala 32:8]
  wire  _GEN_349 = _T_31 ? 1'h0 : _GEN_342; // @[Conditional.scala 39:67 PEArray.scala 208:12]
  wire  _GEN_459 = _T_22 | _GEN_349; // @[Conditional.scala 39:67 PEArray.scala 32:8]
  wire  _GEN_463 = _T_16 ? 1'h0 : _GEN_459; // @[Conditional.scala 39:67]
  wire  _GEN_572 = _T_12 | _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 149:12]
  wire  sel1 = _T_3 | _GEN_572; // @[Conditional.scala 40:58 PEArray.scala 108:12]
  wire [15:0] MAC_out = FP16MAC_io_out; // @[PEArray.scala 47:21 PEArray.scala 85:11]
  wire  _GEN_465 = _T_16 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 177:12]
  wire  _GEN_580 = _T_12 | _GEN_465; // @[Conditional.scala 39:67 PEArray.scala 34:8]
  wire  sel3 = _T_3 | _GEN_580; // @[Conditional.scala 40:58 PEArray.scala 110:12]
  wire [1:0] _GEN_344 = _T_41 ? 2'h2 : 2'h0; // @[Conditional.scala 39:67 PEArray.scala 233:12 PEArray.scala 35:8]
  wire [1:0] _GEN_351 = _T_31 ? 2'h2 : _GEN_344; // @[Conditional.scala 39:67 PEArray.scala 210:12]
  wire [1:0] _GEN_461 = _T_22 ? 2'h0 : _GEN_351; // @[Conditional.scala 39:67 PEArray.scala 35:8]
  wire [1:0] _GEN_466 = _T_16 ? 2'h0 : _GEN_461; // @[Conditional.scala 39:67 PEArray.scala 178:12]
  wire [1:0] _GEN_574 = _T_12 ? 2'h1 : _GEN_466; // @[Conditional.scala 39:67]
  wire [1:0] sel4 = _T_3 ? 2'h0 : _GEN_574; // @[Conditional.scala 40:58 PEArray.scala 111:12]
  wire [15:0] _GEN_3 = sel4 == 2'h2 ? io_FromL1 : 16'h0; // @[PEArray.scala 65:28 PEArray.scala 66:15 PEArray.scala 69:15]
  wire [15:0] _GEN_4 = sel4 == 2'h1 ? io_FromAbovePE : _GEN_3; // @[PEArray.scala 62:28 PEArray.scala 63:15]
  wire [15:0] mux4out = sel4 == 2'h0 ? 16'h0 : _GEN_4; // @[PEArray.scala 59:22 PEArray.scala 60:13]
  wire [15:0] _GEN_7 = 6'h1 == L0Index ? L0Memory_1 : L0Memory_0; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_8 = 6'h2 == L0Index ? L0Memory_2 : _GEN_7; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_9 = 6'h3 == L0Index ? L0Memory_3 : _GEN_8; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_10 = 6'h4 == L0Index ? L0Memory_4 : _GEN_9; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_11 = 6'h5 == L0Index ? L0Memory_5 : _GEN_10; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_12 = 6'h6 == L0Index ? L0Memory_6 : _GEN_11; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_13 = 6'h7 == L0Index ? L0Memory_7 : _GEN_12; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_14 = 6'h8 == L0Index ? L0Memory_8 : _GEN_13; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_15 = 6'h9 == L0Index ? L0Memory_9 : _GEN_14; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_16 = 6'ha == L0Index ? L0Memory_10 : _GEN_15; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_17 = 6'hb == L0Index ? L0Memory_11 : _GEN_16; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_18 = 6'hc == L0Index ? L0Memory_12 : _GEN_17; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_19 = 6'hd == L0Index ? L0Memory_13 : _GEN_18; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_20 = 6'he == L0Index ? L0Memory_14 : _GEN_19; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_21 = 6'hf == L0Index ? L0Memory_15 : _GEN_20; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_22 = 6'h10 == L0Index ? L0Memory_16 : _GEN_21; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_23 = 6'h11 == L0Index ? L0Memory_17 : _GEN_22; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_24 = 6'h12 == L0Index ? L0Memory_18 : _GEN_23; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_25 = 6'h13 == L0Index ? L0Memory_19 : _GEN_24; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_26 = 6'h14 == L0Index ? L0Memory_20 : _GEN_25; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_27 = 6'h15 == L0Index ? L0Memory_21 : _GEN_26; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_28 = 6'h16 == L0Index ? L0Memory_22 : _GEN_27; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_29 = 6'h17 == L0Index ? L0Memory_23 : _GEN_28; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_30 = 6'h18 == L0Index ? L0Memory_24 : _GEN_29; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_31 = 6'h19 == L0Index ? L0Memory_25 : _GEN_30; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_32 = 6'h1a == L0Index ? L0Memory_26 : _GEN_31; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_33 = 6'h1b == L0Index ? L0Memory_27 : _GEN_32; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_34 = 6'h1c == L0Index ? L0Memory_28 : _GEN_33; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_35 = 6'h1d == L0Index ? L0Memory_29 : _GEN_34; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_36 = 6'h1e == L0Index ? L0Memory_30 : _GEN_35; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_37 = 6'h1f == L0Index ? L0Memory_31 : _GEN_36; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_38 = 6'h20 == L0Index ? L0Memory_32 : _GEN_37; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_39 = 6'h21 == L0Index ? L0Memory_33 : _GEN_38; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_40 = 6'h22 == L0Index ? L0Memory_34 : _GEN_39; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_41 = 6'h23 == L0Index ? L0Memory_35 : _GEN_40; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_42 = 6'h24 == L0Index ? L0Memory_36 : _GEN_41; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_43 = 6'h25 == L0Index ? L0Memory_37 : _GEN_42; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_44 = 6'h26 == L0Index ? L0Memory_38 : _GEN_43; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_45 = 6'h27 == L0Index ? L0Memory_39 : _GEN_44; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_46 = 6'h28 == L0Index ? L0Memory_40 : _GEN_45; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_47 = 6'h29 == L0Index ? L0Memory_41 : _GEN_46; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_48 = 6'h2a == L0Index ? L0Memory_42 : _GEN_47; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_49 = 6'h2b == L0Index ? L0Memory_43 : _GEN_48; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_50 = 6'h2c == L0Index ? L0Memory_44 : _GEN_49; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_51 = 6'h2d == L0Index ? L0Memory_45 : _GEN_50; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_52 = 6'h2e == L0Index ? L0Memory_46 : _GEN_51; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_53 = 6'h2f == L0Index ? L0Memory_47 : _GEN_52; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_54 = 6'h30 == L0Index ? L0Memory_48 : _GEN_53; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_55 = 6'h31 == L0Index ? L0Memory_49 : _GEN_54; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_56 = 6'h32 == L0Index ? L0Memory_50 : _GEN_55; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_57 = 6'h33 == L0Index ? L0Memory_51 : _GEN_56; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_58 = 6'h34 == L0Index ? L0Memory_52 : _GEN_57; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_59 = 6'h35 == L0Index ? L0Memory_53 : _GEN_58; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_60 = 6'h36 == L0Index ? L0Memory_54 : _GEN_59; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_61 = 6'h37 == L0Index ? L0Memory_55 : _GEN_60; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_62 = 6'h38 == L0Index ? L0Memory_56 : _GEN_61; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_63 = 6'h39 == L0Index ? L0Memory_57 : _GEN_62; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_64 = 6'h3a == L0Index ? L0Memory_58 : _GEN_63; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_65 = 6'h3b == L0Index ? L0Memory_59 : _GEN_64; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_66 = 6'h3c == L0Index ? L0Memory_60 : _GEN_65; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_67 = 6'h3d == L0Index ? L0Memory_61 : _GEN_66; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_68 = 6'h3e == L0Index ? L0Memory_62 : _GEN_67; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_69 = 6'h3f == L0Index ? L0Memory_63 : _GEN_68; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [6:0] _GEN_793 = {{1'd0}, L0Index}; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_70 = 7'h40 == _GEN_793 ? L0Memory_64 : _GEN_69; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_71 = 7'h41 == _GEN_793 ? L0Memory_65 : _GEN_70; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_72 = 7'h42 == _GEN_793 ? L0Memory_66 : _GEN_71; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_73 = 7'h43 == _GEN_793 ? L0Memory_67 : _GEN_72; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_74 = 7'h44 == _GEN_793 ? L0Memory_68 : _GEN_73; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_75 = 7'h45 == _GEN_793 ? L0Memory_69 : _GEN_74; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_76 = 7'h46 == _GEN_793 ? L0Memory_70 : _GEN_75; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_77 = 7'h47 == _GEN_793 ? L0Memory_71 : _GEN_76; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_78 = 7'h48 == _GEN_793 ? L0Memory_72 : _GEN_77; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_79 = 7'h49 == _GEN_793 ? L0Memory_73 : _GEN_78; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_80 = 7'h4a == _GEN_793 ? L0Memory_74 : _GEN_79; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_81 = 7'h4b == _GEN_793 ? L0Memory_75 : _GEN_80; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_82 = 7'h4c == _GEN_793 ? L0Memory_76 : _GEN_81; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_83 = 7'h4d == _GEN_793 ? L0Memory_77 : _GEN_82; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_84 = 7'h4e == _GEN_793 ? L0Memory_78 : _GEN_83; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_85 = 7'h4f == _GEN_793 ? L0Memory_79 : _GEN_84; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_86 = 7'h50 == _GEN_793 ? L0Memory_80 : _GEN_85; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_87 = 7'h51 == _GEN_793 ? L0Memory_81 : _GEN_86; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_88 = 7'h52 == _GEN_793 ? L0Memory_82 : _GEN_87; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_89 = 7'h53 == _GEN_793 ? L0Memory_83 : _GEN_88; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_90 = 7'h54 == _GEN_793 ? L0Memory_84 : _GEN_89; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_91 = 7'h55 == _GEN_793 ? L0Memory_85 : _GEN_90; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_92 = 7'h56 == _GEN_793 ? L0Memory_86 : _GEN_91; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_93 = 7'h57 == _GEN_793 ? L0Memory_87 : _GEN_92; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_94 = 7'h58 == _GEN_793 ? L0Memory_88 : _GEN_93; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_95 = 7'h59 == _GEN_793 ? L0Memory_89 : _GEN_94; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_96 = 7'h5a == _GEN_793 ? L0Memory_90 : _GEN_95; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_97 = 7'h5b == _GEN_793 ? L0Memory_91 : _GEN_96; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_98 = 7'h5c == _GEN_793 ? L0Memory_92 : _GEN_97; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_99 = 7'h5d == _GEN_793 ? L0Memory_93 : _GEN_98; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_100 = 7'h5e == _GEN_793 ? L0Memory_94 : _GEN_99; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_101 = 7'h5f == _GEN_793 ? L0Memory_95 : _GEN_100; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_102 = 7'h60 == _GEN_793 ? L0Memory_96 : _GEN_101; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_103 = 7'h61 == _GEN_793 ? L0Memory_97 : _GEN_102; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_104 = 7'h62 == _GEN_793 ? L0Memory_98 : _GEN_103; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_105 = 7'h63 == _GEN_793 ? L0Memory_99 : _GEN_104; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire  _GEN_575 = _T_12 ? 1'h0 : _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 157:12]
  wire  sel5 = _T_3 ? 1'h0 : _GEN_575; // @[Conditional.scala 40:58 PEArray.scala 112:12]
  reg [15:0] mux2out_reg; // @[PEArray.scala 90:28]
  reg [15:0] mux3out_reg; // @[PEArray.scala 91:28]
  reg [9:0] count; // @[PEArray.scala 101:22]
  reg [9:0] count_max; // @[PEArray.scala 102:22]
  reg [5:0] L0index_begin; // @[PEArray.scala 103:26]
  reg [5:0] GRU_out_width; // @[PEArray.scala 104:26]
  wire  _T_6 = 3'h0 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_7 = 3'h1 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_8 = 3'h2 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_9 = 3'h3 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_10 = 3'h4 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_11 = 3'h5 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_109 = _T_11 ? 3'h5 : state; // @[Conditional.scala 39:67 PEArray.scala 140:19 PEArray.scala 100:22]
  wire [2:0] _GEN_110 = _T_10 ? 3'h4 : _GEN_109; // @[Conditional.scala 39:67 PEArray.scala 136:19]
  wire [2:0] _GEN_111 = _T_9 ? 3'h3 : _GEN_110; // @[Conditional.scala 39:67 PEArray.scala 132:19]
  wire [2:0] _GEN_112 = _T_8 ? 3'h2 : _GEN_111; // @[Conditional.scala 39:67 PEArray.scala 128:19]
  wire [2:0] _GEN_113 = _T_7 ? 3'h1 : _GEN_112; // @[Conditional.scala 39:67 PEArray.scala 124:19]
  wire [7:0] _GEN_118 = io_control_signal_mask[2] ? io_control_signal_gru_out_width : {{2'd0}, GRU_out_width}; // @[PEArray.scala 116:57 PEArray.scala 145:23 PEArray.scala 104:26]
  wire [9:0] _count_T_1 = count + 10'h1; // @[PEArray.scala 162:24]
  wire [9:0] _GEN_120 = count != 10'h33 ? _count_T_1 : count; // @[PEArray.scala 161:27 PEArray.scala 162:15 PEArray.scala 101:22]
  wire [9:0] _GEN_124 = count != 10'h188 ? _count_T_1 : count; // @[PEArray.scala 183:28 PEArray.scala 184:15 PEArray.scala 101:22]
  wire [9:0] _GEN_125 = count == 10'h188 ? 10'h0 : _GEN_124; // @[PEArray.scala 186:28 PEArray.scala 187:15]
  wire [2:0] _GEN_126 = count == 10'h188 ? 3'h0 : state; // @[PEArray.scala 186:28 PEArray.scala 188:15 PEArray.scala 100:22]
  wire [9:0] _GEN_127 = count != count_max ? _count_T_1 : count; // @[PEArray.scala 192:32 PEArray.scala 193:15 PEArray.scala 101:22]
  wire [5:0] _GEN_128 = count == 10'h0 ? L0index_begin : L0Index; // @[PEArray.scala 195:26 PEArray.scala 196:17 PEArray.scala 39:24]
  wire [9:0] _T_27 = count_max - 10'h1; // @[PEArray.scala 198:51]
  wire [15:0] _GEN_129 = 6'h0 == L0Index ? io_FromL1 : L0Memory_0; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_130 = 6'h1 == L0Index ? io_FromL1 : L0Memory_1; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_131 = 6'h2 == L0Index ? io_FromL1 : L0Memory_2; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_132 = 6'h3 == L0Index ? io_FromL1 : L0Memory_3; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_133 = 6'h4 == L0Index ? io_FromL1 : L0Memory_4; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_134 = 6'h5 == L0Index ? io_FromL1 : L0Memory_5; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_135 = 6'h6 == L0Index ? io_FromL1 : L0Memory_6; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_136 = 6'h7 == L0Index ? io_FromL1 : L0Memory_7; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_137 = 6'h8 == L0Index ? io_FromL1 : L0Memory_8; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_138 = 6'h9 == L0Index ? io_FromL1 : L0Memory_9; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_139 = 6'ha == L0Index ? io_FromL1 : L0Memory_10; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_140 = 6'hb == L0Index ? io_FromL1 : L0Memory_11; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_141 = 6'hc == L0Index ? io_FromL1 : L0Memory_12; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_142 = 6'hd == L0Index ? io_FromL1 : L0Memory_13; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_143 = 6'he == L0Index ? io_FromL1 : L0Memory_14; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_144 = 6'hf == L0Index ? io_FromL1 : L0Memory_15; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_145 = 6'h10 == L0Index ? io_FromL1 : L0Memory_16; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_146 = 6'h11 == L0Index ? io_FromL1 : L0Memory_17; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_147 = 6'h12 == L0Index ? io_FromL1 : L0Memory_18; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_148 = 6'h13 == L0Index ? io_FromL1 : L0Memory_19; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_149 = 6'h14 == L0Index ? io_FromL1 : L0Memory_20; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_150 = 6'h15 == L0Index ? io_FromL1 : L0Memory_21; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_151 = 6'h16 == L0Index ? io_FromL1 : L0Memory_22; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_152 = 6'h17 == L0Index ? io_FromL1 : L0Memory_23; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_153 = 6'h18 == L0Index ? io_FromL1 : L0Memory_24; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_154 = 6'h19 == L0Index ? io_FromL1 : L0Memory_25; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_155 = 6'h1a == L0Index ? io_FromL1 : L0Memory_26; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_156 = 6'h1b == L0Index ? io_FromL1 : L0Memory_27; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_157 = 6'h1c == L0Index ? io_FromL1 : L0Memory_28; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_158 = 6'h1d == L0Index ? io_FromL1 : L0Memory_29; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_159 = 6'h1e == L0Index ? io_FromL1 : L0Memory_30; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_160 = 6'h1f == L0Index ? io_FromL1 : L0Memory_31; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_161 = 6'h20 == L0Index ? io_FromL1 : L0Memory_32; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_162 = 6'h21 == L0Index ? io_FromL1 : L0Memory_33; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_163 = 6'h22 == L0Index ? io_FromL1 : L0Memory_34; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_164 = 6'h23 == L0Index ? io_FromL1 : L0Memory_35; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_165 = 6'h24 == L0Index ? io_FromL1 : L0Memory_36; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_166 = 6'h25 == L0Index ? io_FromL1 : L0Memory_37; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_167 = 6'h26 == L0Index ? io_FromL1 : L0Memory_38; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_168 = 6'h27 == L0Index ? io_FromL1 : L0Memory_39; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_169 = 6'h28 == L0Index ? io_FromL1 : L0Memory_40; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_170 = 6'h29 == L0Index ? io_FromL1 : L0Memory_41; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_171 = 6'h2a == L0Index ? io_FromL1 : L0Memory_42; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_172 = 6'h2b == L0Index ? io_FromL1 : L0Memory_43; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_173 = 6'h2c == L0Index ? io_FromL1 : L0Memory_44; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_174 = 6'h2d == L0Index ? io_FromL1 : L0Memory_45; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_175 = 6'h2e == L0Index ? io_FromL1 : L0Memory_46; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_176 = 6'h2f == L0Index ? io_FromL1 : L0Memory_47; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_177 = 6'h30 == L0Index ? io_FromL1 : L0Memory_48; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_178 = 6'h31 == L0Index ? io_FromL1 : L0Memory_49; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_179 = 6'h32 == L0Index ? io_FromL1 : L0Memory_50; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_180 = 6'h33 == L0Index ? io_FromL1 : L0Memory_51; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_181 = 6'h34 == L0Index ? io_FromL1 : L0Memory_52; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_182 = 6'h35 == L0Index ? io_FromL1 : L0Memory_53; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_183 = 6'h36 == L0Index ? io_FromL1 : L0Memory_54; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_184 = 6'h37 == L0Index ? io_FromL1 : L0Memory_55; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_185 = 6'h38 == L0Index ? io_FromL1 : L0Memory_56; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_186 = 6'h39 == L0Index ? io_FromL1 : L0Memory_57; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_187 = 6'h3a == L0Index ? io_FromL1 : L0Memory_58; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_188 = 6'h3b == L0Index ? io_FromL1 : L0Memory_59; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_189 = 6'h3c == L0Index ? io_FromL1 : L0Memory_60; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_190 = 6'h3d == L0Index ? io_FromL1 : L0Memory_61; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_191 = 6'h3e == L0Index ? io_FromL1 : L0Memory_62; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_192 = 6'h3f == L0Index ? io_FromL1 : L0Memory_63; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_193 = 7'h40 == _GEN_793 ? io_FromL1 : L0Memory_64; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_194 = 7'h41 == _GEN_793 ? io_FromL1 : L0Memory_65; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_195 = 7'h42 == _GEN_793 ? io_FromL1 : L0Memory_66; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_196 = 7'h43 == _GEN_793 ? io_FromL1 : L0Memory_67; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_197 = 7'h44 == _GEN_793 ? io_FromL1 : L0Memory_68; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_198 = 7'h45 == _GEN_793 ? io_FromL1 : L0Memory_69; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_199 = 7'h46 == _GEN_793 ? io_FromL1 : L0Memory_70; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_200 = 7'h47 == _GEN_793 ? io_FromL1 : L0Memory_71; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_201 = 7'h48 == _GEN_793 ? io_FromL1 : L0Memory_72; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_202 = 7'h49 == _GEN_793 ? io_FromL1 : L0Memory_73; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_203 = 7'h4a == _GEN_793 ? io_FromL1 : L0Memory_74; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_204 = 7'h4b == _GEN_793 ? io_FromL1 : L0Memory_75; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_205 = 7'h4c == _GEN_793 ? io_FromL1 : L0Memory_76; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_206 = 7'h4d == _GEN_793 ? io_FromL1 : L0Memory_77; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_207 = 7'h4e == _GEN_793 ? io_FromL1 : L0Memory_78; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_208 = 7'h4f == _GEN_793 ? io_FromL1 : L0Memory_79; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_209 = 7'h50 == _GEN_793 ? io_FromL1 : L0Memory_80; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_210 = 7'h51 == _GEN_793 ? io_FromL1 : L0Memory_81; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_211 = 7'h52 == _GEN_793 ? io_FromL1 : L0Memory_82; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_212 = 7'h53 == _GEN_793 ? io_FromL1 : L0Memory_83; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_213 = 7'h54 == _GEN_793 ? io_FromL1 : L0Memory_84; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_214 = 7'h55 == _GEN_793 ? io_FromL1 : L0Memory_85; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_215 = 7'h56 == _GEN_793 ? io_FromL1 : L0Memory_86; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_216 = 7'h57 == _GEN_793 ? io_FromL1 : L0Memory_87; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_217 = 7'h58 == _GEN_793 ? io_FromL1 : L0Memory_88; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_218 = 7'h59 == _GEN_793 ? io_FromL1 : L0Memory_89; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_219 = 7'h5a == _GEN_793 ? io_FromL1 : L0Memory_90; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_220 = 7'h5b == _GEN_793 ? io_FromL1 : L0Memory_91; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_221 = 7'h5c == _GEN_793 ? io_FromL1 : L0Memory_92; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_222 = 7'h5d == _GEN_793 ? io_FromL1 : L0Memory_93; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_223 = 7'h5e == _GEN_793 ? io_FromL1 : L0Memory_94; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_224 = 7'h5f == _GEN_793 ? io_FromL1 : L0Memory_95; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_225 = 7'h60 == _GEN_793 ? io_FromL1 : L0Memory_96; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_226 = 7'h61 == _GEN_793 ? io_FromL1 : L0Memory_97; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_227 = 7'h62 == _GEN_793 ? io_FromL1 : L0Memory_98; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_228 = 7'h63 == _GEN_793 ? io_FromL1 : L0Memory_99; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [5:0] _L0Index_T_2 = L0Index + 6'h1; // @[PEArray.scala 200:28]
  wire [15:0] _GEN_229 = count >= 10'h1 & count <= _T_27 ? _GEN_129 : L0Memory_0; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_230 = count >= 10'h1 & count <= _T_27 ? _GEN_130 : L0Memory_1; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_231 = count >= 10'h1 & count <= _T_27 ? _GEN_131 : L0Memory_2; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_232 = count >= 10'h1 & count <= _T_27 ? _GEN_132 : L0Memory_3; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_233 = count >= 10'h1 & count <= _T_27 ? _GEN_133 : L0Memory_4; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_234 = count >= 10'h1 & count <= _T_27 ? _GEN_134 : L0Memory_5; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_235 = count >= 10'h1 & count <= _T_27 ? _GEN_135 : L0Memory_6; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_236 = count >= 10'h1 & count <= _T_27 ? _GEN_136 : L0Memory_7; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_237 = count >= 10'h1 & count <= _T_27 ? _GEN_137 : L0Memory_8; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_238 = count >= 10'h1 & count <= _T_27 ? _GEN_138 : L0Memory_9; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_239 = count >= 10'h1 & count <= _T_27 ? _GEN_139 : L0Memory_10; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_240 = count >= 10'h1 & count <= _T_27 ? _GEN_140 : L0Memory_11; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_241 = count >= 10'h1 & count <= _T_27 ? _GEN_141 : L0Memory_12; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_242 = count >= 10'h1 & count <= _T_27 ? _GEN_142 : L0Memory_13; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_243 = count >= 10'h1 & count <= _T_27 ? _GEN_143 : L0Memory_14; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_244 = count >= 10'h1 & count <= _T_27 ? _GEN_144 : L0Memory_15; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_245 = count >= 10'h1 & count <= _T_27 ? _GEN_145 : L0Memory_16; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_246 = count >= 10'h1 & count <= _T_27 ? _GEN_146 : L0Memory_17; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_247 = count >= 10'h1 & count <= _T_27 ? _GEN_147 : L0Memory_18; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_248 = count >= 10'h1 & count <= _T_27 ? _GEN_148 : L0Memory_19; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_249 = count >= 10'h1 & count <= _T_27 ? _GEN_149 : L0Memory_20; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_250 = count >= 10'h1 & count <= _T_27 ? _GEN_150 : L0Memory_21; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_251 = count >= 10'h1 & count <= _T_27 ? _GEN_151 : L0Memory_22; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_252 = count >= 10'h1 & count <= _T_27 ? _GEN_152 : L0Memory_23; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_253 = count >= 10'h1 & count <= _T_27 ? _GEN_153 : L0Memory_24; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_254 = count >= 10'h1 & count <= _T_27 ? _GEN_154 : L0Memory_25; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_255 = count >= 10'h1 & count <= _T_27 ? _GEN_155 : L0Memory_26; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_256 = count >= 10'h1 & count <= _T_27 ? _GEN_156 : L0Memory_27; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_257 = count >= 10'h1 & count <= _T_27 ? _GEN_157 : L0Memory_28; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_258 = count >= 10'h1 & count <= _T_27 ? _GEN_158 : L0Memory_29; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_259 = count >= 10'h1 & count <= _T_27 ? _GEN_159 : L0Memory_30; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_260 = count >= 10'h1 & count <= _T_27 ? _GEN_160 : L0Memory_31; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_261 = count >= 10'h1 & count <= _T_27 ? _GEN_161 : L0Memory_32; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_262 = count >= 10'h1 & count <= _T_27 ? _GEN_162 : L0Memory_33; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_263 = count >= 10'h1 & count <= _T_27 ? _GEN_163 : L0Memory_34; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_264 = count >= 10'h1 & count <= _T_27 ? _GEN_164 : L0Memory_35; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_265 = count >= 10'h1 & count <= _T_27 ? _GEN_165 : L0Memory_36; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_266 = count >= 10'h1 & count <= _T_27 ? _GEN_166 : L0Memory_37; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_267 = count >= 10'h1 & count <= _T_27 ? _GEN_167 : L0Memory_38; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_268 = count >= 10'h1 & count <= _T_27 ? _GEN_168 : L0Memory_39; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_269 = count >= 10'h1 & count <= _T_27 ? _GEN_169 : L0Memory_40; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_270 = count >= 10'h1 & count <= _T_27 ? _GEN_170 : L0Memory_41; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_271 = count >= 10'h1 & count <= _T_27 ? _GEN_171 : L0Memory_42; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_272 = count >= 10'h1 & count <= _T_27 ? _GEN_172 : L0Memory_43; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_273 = count >= 10'h1 & count <= _T_27 ? _GEN_173 : L0Memory_44; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_274 = count >= 10'h1 & count <= _T_27 ? _GEN_174 : L0Memory_45; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_275 = count >= 10'h1 & count <= _T_27 ? _GEN_175 : L0Memory_46; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_276 = count >= 10'h1 & count <= _T_27 ? _GEN_176 : L0Memory_47; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_277 = count >= 10'h1 & count <= _T_27 ? _GEN_177 : L0Memory_48; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_278 = count >= 10'h1 & count <= _T_27 ? _GEN_178 : L0Memory_49; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_279 = count >= 10'h1 & count <= _T_27 ? _GEN_179 : L0Memory_50; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_280 = count >= 10'h1 & count <= _T_27 ? _GEN_180 : L0Memory_51; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_281 = count >= 10'h1 & count <= _T_27 ? _GEN_181 : L0Memory_52; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_282 = count >= 10'h1 & count <= _T_27 ? _GEN_182 : L0Memory_53; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_283 = count >= 10'h1 & count <= _T_27 ? _GEN_183 : L0Memory_54; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_284 = count >= 10'h1 & count <= _T_27 ? _GEN_184 : L0Memory_55; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_285 = count >= 10'h1 & count <= _T_27 ? _GEN_185 : L0Memory_56; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_286 = count >= 10'h1 & count <= _T_27 ? _GEN_186 : L0Memory_57; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_287 = count >= 10'h1 & count <= _T_27 ? _GEN_187 : L0Memory_58; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_288 = count >= 10'h1 & count <= _T_27 ? _GEN_188 : L0Memory_59; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_289 = count >= 10'h1 & count <= _T_27 ? _GEN_189 : L0Memory_60; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_290 = count >= 10'h1 & count <= _T_27 ? _GEN_190 : L0Memory_61; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_291 = count >= 10'h1 & count <= _T_27 ? _GEN_191 : L0Memory_62; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_292 = count >= 10'h1 & count <= _T_27 ? _GEN_192 : L0Memory_63; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_293 = count >= 10'h1 & count <= _T_27 ? _GEN_193 : L0Memory_64; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_294 = count >= 10'h1 & count <= _T_27 ? _GEN_194 : L0Memory_65; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_295 = count >= 10'h1 & count <= _T_27 ? _GEN_195 : L0Memory_66; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_296 = count >= 10'h1 & count <= _T_27 ? _GEN_196 : L0Memory_67; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_297 = count >= 10'h1 & count <= _T_27 ? _GEN_197 : L0Memory_68; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_298 = count >= 10'h1 & count <= _T_27 ? _GEN_198 : L0Memory_69; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_299 = count >= 10'h1 & count <= _T_27 ? _GEN_199 : L0Memory_70; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_300 = count >= 10'h1 & count <= _T_27 ? _GEN_200 : L0Memory_71; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_301 = count >= 10'h1 & count <= _T_27 ? _GEN_201 : L0Memory_72; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_302 = count >= 10'h1 & count <= _T_27 ? _GEN_202 : L0Memory_73; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_303 = count >= 10'h1 & count <= _T_27 ? _GEN_203 : L0Memory_74; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_304 = count >= 10'h1 & count <= _T_27 ? _GEN_204 : L0Memory_75; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_305 = count >= 10'h1 & count <= _T_27 ? _GEN_205 : L0Memory_76; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_306 = count >= 10'h1 & count <= _T_27 ? _GEN_206 : L0Memory_77; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_307 = count >= 10'h1 & count <= _T_27 ? _GEN_207 : L0Memory_78; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_308 = count >= 10'h1 & count <= _T_27 ? _GEN_208 : L0Memory_79; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_309 = count >= 10'h1 & count <= _T_27 ? _GEN_209 : L0Memory_80; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_310 = count >= 10'h1 & count <= _T_27 ? _GEN_210 : L0Memory_81; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_311 = count >= 10'h1 & count <= _T_27 ? _GEN_211 : L0Memory_82; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_312 = count >= 10'h1 & count <= _T_27 ? _GEN_212 : L0Memory_83; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_313 = count >= 10'h1 & count <= _T_27 ? _GEN_213 : L0Memory_84; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_314 = count >= 10'h1 & count <= _T_27 ? _GEN_214 : L0Memory_85; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_315 = count >= 10'h1 & count <= _T_27 ? _GEN_215 : L0Memory_86; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_316 = count >= 10'h1 & count <= _T_27 ? _GEN_216 : L0Memory_87; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_317 = count >= 10'h1 & count <= _T_27 ? _GEN_217 : L0Memory_88; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_318 = count >= 10'h1 & count <= _T_27 ? _GEN_218 : L0Memory_89; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_319 = count >= 10'h1 & count <= _T_27 ? _GEN_219 : L0Memory_90; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_320 = count >= 10'h1 & count <= _T_27 ? _GEN_220 : L0Memory_91; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_321 = count >= 10'h1 & count <= _T_27 ? _GEN_221 : L0Memory_92; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_322 = count >= 10'h1 & count <= _T_27 ? _GEN_222 : L0Memory_93; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_323 = count >= 10'h1 & count <= _T_27 ? _GEN_223 : L0Memory_94; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_324 = count >= 10'h1 & count <= _T_27 ? _GEN_224 : L0Memory_95; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_325 = count >= 10'h1 & count <= _T_27 ? _GEN_225 : L0Memory_96; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_326 = count >= 10'h1 & count <= _T_27 ? _GEN_226 : L0Memory_97; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_327 = count >= 10'h1 & count <= _T_27 ? _GEN_227 : L0Memory_98; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_328 = count >= 10'h1 & count <= _T_27 ? _GEN_228 : L0Memory_99; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [5:0] _GEN_329 = count >= 10'h1 & count <= _T_27 ? _L0Index_T_2 : _GEN_128; // @[PEArray.scala 198:59 PEArray.scala 200:17]
  wire [9:0] _GEN_330 = count == count_max ? 10'h0 : _GEN_127; // @[PEArray.scala 202:32 PEArray.scala 203:15]
  wire [2:0] _GEN_331 = count == count_max ? 3'h0 : state; // @[PEArray.scala 202:32 PEArray.scala 204:15 PEArray.scala 100:22]
  wire [9:0] _GEN_865 = {{4'd0}, GRU_out_width}; // @[PEArray.scala 220:19]
  wire [9:0] _GEN_0 = count % _GEN_865; // @[PEArray.scala 220:19]
  wire [5:0] _T_36 = _GEN_0[5:0]; // @[PEArray.scala 220:19]
  wire [5:0] _T_38 = GRU_out_width - 6'h1; // @[PEArray.scala 220:55]
  wire [5:0] _GEN_334 = _T_36 == _T_38 ? _L0Index_T_2 : L0index_begin; // @[PEArray.scala 220:62 PEArray.scala 221:17 PEArray.scala 214:15]
  wire [5:0] _GEN_346 = _T_41 ? _GEN_334 : L0Index; // @[Conditional.scala 39:67 PEArray.scala 39:24]
  wire [9:0] _GEN_347 = _T_41 ? _GEN_330 : count; // @[Conditional.scala 39:67 PEArray.scala 101:22]
  wire [2:0] _GEN_348 = _T_41 ? _GEN_331 : state; // @[Conditional.scala 39:67 PEArray.scala 100:22]
  wire [5:0] _GEN_353 = _T_31 ? _GEN_334 : _GEN_346; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_354 = _T_31 ? _GEN_330 : _GEN_347; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_355 = _T_31 ? _GEN_331 : _GEN_348; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_356 = _T_22 ? _GEN_330 : _GEN_354; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_357 = _T_22 ? _GEN_329 : _GEN_353; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_458 = _T_22 ? _GEN_331 : _GEN_355; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_690 = _T_3 ? _GEN_118 : {{2'd0}, GRU_out_width}; // @[Conditional.scala 40:58 PEArray.scala 104:26]
  FP16MulAdder FP16MAC ( // @[PEArray.scala 72:23]
    .io_a(FP16MAC_io_a),
    .io_b(FP16MAC_io_b),
    .io_c(FP16MAC_io_c),
    .io_out(FP16MAC_io_out)
  );
  assign io_ToRightPE = mux3out_reg; // @[PEArray.scala 95:16]
  assign io_ToBelowPE = mux2out_reg; // @[PEArray.scala 94:16]
  assign FP16MAC_io_a = sel1 ? io_FromL1 : io_FromLeftPE; // @[PEArray.scala 50:14 PEArray.scala 50:23 PEArray.scala 51:24]
  assign FP16MAC_io_b = sel5 ? mux4out : _GEN_105; // @[PEArray.scala 77:13 PEArray.scala 78:18 PEArray.scala 81:18]
  assign FP16MAC_io_c = sel5 ? _GEN_105 : mux4out; // @[PEArray.scala 77:13 PEArray.scala 79:18 PEArray.scala 82:18]
  always @(posedge clock) begin
    if (reset) begin // @[PEArray.scala 39:24]
      L0Index <= 6'h0; // @[PEArray.scala 39:24]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h2; // @[PEArray.scala 159:15]
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        L0Index <= 6'hc; // @[PEArray.scala 181:15]
      end else begin
        L0Index <= _GEN_357;
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_0 <= _GEN_229;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_1 <= _GEN_230;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_2 <= _GEN_231;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_3 <= _GEN_232;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_4 <= _GEN_233;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_5 <= _GEN_234;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_6 <= _GEN_235;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_7 <= _GEN_236;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_8 <= _GEN_237;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_9 <= _GEN_238;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_10 <= _GEN_239;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_11 <= _GEN_240;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_12 <= _GEN_241;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_13 <= _GEN_242;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_14 <= _GEN_243;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_15 <= _GEN_244;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_16 <= _GEN_245;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_17 <= _GEN_246;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_18 <= _GEN_247;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_19 <= _GEN_248;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_20 <= _GEN_249;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_21 <= _GEN_250;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_22 <= _GEN_251;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_23 <= _GEN_252;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_24 <= _GEN_253;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_25 <= _GEN_254;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_26 <= _GEN_255;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_27 <= _GEN_256;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_28 <= _GEN_257;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_29 <= _GEN_258;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_30 <= _GEN_259;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_31 <= _GEN_260;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_32 <= _GEN_261;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_33 <= _GEN_262;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_34 <= _GEN_263;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_35 <= _GEN_264;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_36 <= _GEN_265;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_37 <= _GEN_266;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_38 <= _GEN_267;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_39 <= _GEN_268;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_40 <= _GEN_269;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_41 <= _GEN_270;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_42 <= _GEN_271;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_43 <= _GEN_272;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_44 <= _GEN_273;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_45 <= _GEN_274;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_46 <= _GEN_275;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_47 <= _GEN_276;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_48 <= _GEN_277;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_49 <= _GEN_278;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_50 <= _GEN_279;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_51 <= _GEN_280;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_52 <= _GEN_281;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_53 <= _GEN_282;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_54 <= _GEN_283;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_55 <= _GEN_284;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_56 <= _GEN_285;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_57 <= _GEN_286;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_58 <= _GEN_287;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_59 <= _GEN_288;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_60 <= _GEN_289;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_61 <= _GEN_290;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_62 <= _GEN_291;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_63 <= _GEN_292;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_64 <= _GEN_293;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_65 <= _GEN_294;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_66 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_67 <= _GEN_296;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_68 <= _GEN_297;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_69 <= _GEN_298;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_70 <= _GEN_299;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_71 <= _GEN_300;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_72 <= _GEN_301;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_73 <= _GEN_302;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_74 <= _GEN_303;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_75 <= _GEN_304;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_76 <= _GEN_305;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_77 <= _GEN_306;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_78 <= _GEN_307;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_79 <= _GEN_308;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_80 <= _GEN_309;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_81 <= _GEN_310;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_82 <= _GEN_311;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_83 <= _GEN_312;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_84 <= _GEN_313;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_85 <= _GEN_314;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_86 <= _GEN_315;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_87 <= _GEN_316;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_88 <= _GEN_317;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_89 <= _GEN_318;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_90 <= _GEN_319;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_91 <= _GEN_320;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_92 <= _GEN_321;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_93 <= _GEN_322;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_94 <= _GEN_323;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_95 <= _GEN_324;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_96 <= _GEN_325;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_97 <= _GEN_326;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_98 <= _GEN_327;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_99 <= _GEN_328;
          end
        end
      end
    end
    if (reset) begin // @[PEArray.scala 100:22]
      state <= 3'h0; // @[PEArray.scala 100:22]
    end else if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[2]) begin // @[PEArray.scala 116:57]
        if (_T_6) begin // @[Conditional.scala 40:58]
          state <= 3'h0; // @[PEArray.scala 120:19]
        end else begin
          state <= _GEN_113;
        end
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      if (count == 10'h33) begin // @[PEArray.scala 164:27]
        state <= 3'h0; // @[PEArray.scala 166:15]
      end
    end else if (_T_16) begin // @[Conditional.scala 39:67]
      state <= _GEN_126;
    end else begin
      state <= _GEN_458;
    end
    if (reset) begin // @[PEArray.scala 90:28]
      mux2out_reg <= 16'h0; // @[PEArray.scala 90:28]
    end else begin
      mux2out_reg <= MAC_out; // @[PEArray.scala 90:28]
    end
    if (reset) begin // @[PEArray.scala 91:28]
      mux3out_reg <= 16'h0; // @[PEArray.scala 91:28]
    end else if (sel3) begin // @[PEArray.scala 56:14]
      mux3out_reg <= MAC_out; // @[PEArray.scala 56:23]
    end else if (sel1) begin // @[PEArray.scala 50:14]
      mux3out_reg <= io_FromL1; // @[PEArray.scala 50:23]
    end else begin
      mux3out_reg <= io_FromLeftPE; // @[PEArray.scala 51:24]
    end
    if (reset) begin // @[PEArray.scala 101:22]
      count <= 10'h0; // @[PEArray.scala 101:22]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        if (count == 10'h33) begin // @[PEArray.scala 164:27]
          count <= 10'h0; // @[PEArray.scala 165:15]
        end else begin
          count <= _GEN_120;
        end
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        count <= _GEN_125;
      end else begin
        count <= _GEN_356;
      end
    end
    if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[2]) begin // @[PEArray.scala 116:57]
        count_max <= io_control_signal_count; // @[PEArray.scala 143:19]
      end
    end
    if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[2]) begin // @[PEArray.scala 116:57]
        L0index_begin <= io_control_signal_L0index; // @[PEArray.scala 144:23]
      end
    end
    GRU_out_width <= _GEN_690[5:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  L0Index = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  L0Memory_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  L0Memory_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  L0Memory_2 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  L0Memory_3 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  L0Memory_4 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  L0Memory_5 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  L0Memory_6 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  L0Memory_7 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  L0Memory_8 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  L0Memory_9 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  L0Memory_10 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  L0Memory_11 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  L0Memory_12 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  L0Memory_13 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  L0Memory_14 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  L0Memory_15 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  L0Memory_16 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  L0Memory_17 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  L0Memory_18 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  L0Memory_19 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  L0Memory_20 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  L0Memory_21 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  L0Memory_22 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  L0Memory_23 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  L0Memory_24 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  L0Memory_25 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  L0Memory_26 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  L0Memory_27 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  L0Memory_28 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  L0Memory_29 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  L0Memory_30 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  L0Memory_31 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  L0Memory_32 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  L0Memory_33 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  L0Memory_34 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  L0Memory_35 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  L0Memory_36 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  L0Memory_37 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  L0Memory_38 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  L0Memory_39 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  L0Memory_40 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  L0Memory_41 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  L0Memory_42 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  L0Memory_43 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  L0Memory_44 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  L0Memory_45 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  L0Memory_46 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  L0Memory_47 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  L0Memory_48 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  L0Memory_49 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  L0Memory_50 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  L0Memory_51 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  L0Memory_52 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  L0Memory_53 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  L0Memory_54 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  L0Memory_55 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  L0Memory_56 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  L0Memory_57 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  L0Memory_58 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  L0Memory_59 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  L0Memory_60 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  L0Memory_61 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  L0Memory_62 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  L0Memory_63 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  L0Memory_64 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  L0Memory_65 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  L0Memory_66 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  L0Memory_67 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  L0Memory_68 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  L0Memory_69 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  L0Memory_70 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  L0Memory_71 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  L0Memory_72 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  L0Memory_73 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  L0Memory_74 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  L0Memory_75 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  L0Memory_76 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  L0Memory_77 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  L0Memory_78 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  L0Memory_79 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  L0Memory_80 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  L0Memory_81 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  L0Memory_82 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  L0Memory_83 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  L0Memory_84 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  L0Memory_85 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  L0Memory_86 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  L0Memory_87 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  L0Memory_88 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  L0Memory_89 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  L0Memory_90 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  L0Memory_91 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  L0Memory_92 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  L0Memory_93 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  L0Memory_94 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  L0Memory_95 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  L0Memory_96 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  L0Memory_97 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  L0Memory_98 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  L0Memory_99 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  state = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  mux2out_reg = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  mux3out_reg = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  count = _RAND_104[9:0];
  _RAND_105 = {1{`RANDOM}};
  count_max = _RAND_105[9:0];
  _RAND_106 = {1{`RANDOM}};
  L0index_begin = _RAND_106[5:0];
  _RAND_107 = {1{`RANDOM}};
  GRU_out_width = _RAND_107[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PE_30(
  input         clock,
  input         reset,
  input  [15:0] io_FromAbovePE,
  input  [15:0] io_FromLeftPE,
  input  [15:0] io_FromL1,
  input  [11:0] io_control_signal_mask,
  output [15:0] io_ToRightPE,
  output [15:0] io_ToBelowPE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] FP16MAC_io_a; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_b; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_c; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_out; // @[PEArray.scala 72:23]
  reg [5:0] L0Index; // @[PEArray.scala 39:24]
  reg [15:0] L0Memory_0; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_1; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_2; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_3; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_4; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_5; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_6; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_7; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_8; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_9; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_10; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_11; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_12; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_13; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_14; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_15; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_16; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_17; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_18; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_19; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_20; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_21; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_22; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_23; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_24; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_25; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_26; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_27; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_28; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_29; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_30; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_31; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_32; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_33; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_34; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_35; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_36; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_37; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_38; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_39; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_40; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_41; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_42; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_43; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_44; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_45; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_46; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_47; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_48; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_49; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_50; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_51; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_52; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_53; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_54; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_55; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_56; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_57; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_58; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_59; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_60; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_61; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_62; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_63; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_64; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_65; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_66; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_67; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_68; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_69; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_70; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_71; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_72; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_73; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_74; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_75; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_76; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_77; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_78; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_79; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_80; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_81; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_82; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_83; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_84; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_85; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_86; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_87; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_88; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_89; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_90; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_91; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_92; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_93; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_94; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_95; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_96; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_97; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_98; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_99; // @[PEArray.scala 40:21]
  reg [2:0] state; // @[PEArray.scala 100:22]
  wire  _T_3 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_12 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_16 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_22 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_31 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_41 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_342 = _T_41 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 231:12 PEArray.scala 32:8]
  wire  _GEN_349 = _T_31 ? 1'h0 : _GEN_342; // @[Conditional.scala 39:67 PEArray.scala 208:12]
  wire  _GEN_459 = _T_22 | _GEN_349; // @[Conditional.scala 39:67 PEArray.scala 32:8]
  wire  _GEN_463 = _T_16 ? 1'h0 : _GEN_459; // @[Conditional.scala 39:67]
  wire  _GEN_572 = _T_12 | _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 149:12]
  wire  sel1 = _T_3 | _GEN_572; // @[Conditional.scala 40:58 PEArray.scala 108:12]
  wire [15:0] MAC_out = FP16MAC_io_out; // @[PEArray.scala 47:21 PEArray.scala 85:11]
  wire  _GEN_465 = _T_16 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 177:12]
  wire  _GEN_580 = _T_12 | _GEN_465; // @[Conditional.scala 39:67 PEArray.scala 34:8]
  wire  sel3 = _T_3 | _GEN_580; // @[Conditional.scala 40:58 PEArray.scala 110:12]
  wire [1:0] _GEN_344 = _T_41 ? 2'h2 : 2'h0; // @[Conditional.scala 39:67 PEArray.scala 233:12 PEArray.scala 35:8]
  wire [1:0] _GEN_351 = _T_31 ? 2'h2 : _GEN_344; // @[Conditional.scala 39:67 PEArray.scala 210:12]
  wire [1:0] _GEN_461 = _T_22 ? 2'h0 : _GEN_351; // @[Conditional.scala 39:67 PEArray.scala 35:8]
  wire [1:0] _GEN_466 = _T_16 ? 2'h0 : _GEN_461; // @[Conditional.scala 39:67 PEArray.scala 178:12]
  wire [1:0] _GEN_574 = _T_12 ? 2'h0 : _GEN_466; // @[Conditional.scala 39:67]
  wire [1:0] sel4 = _T_3 ? 2'h0 : _GEN_574; // @[Conditional.scala 40:58 PEArray.scala 111:12]
  wire [15:0] _GEN_3 = sel4 == 2'h2 ? io_FromL1 : 16'h0; // @[PEArray.scala 65:28 PEArray.scala 66:15 PEArray.scala 69:15]
  wire [15:0] _GEN_4 = sel4 == 2'h1 ? io_FromAbovePE : _GEN_3; // @[PEArray.scala 62:28 PEArray.scala 63:15]
  wire [15:0] mux4out = sel4 == 2'h0 ? 16'h0 : _GEN_4; // @[PEArray.scala 59:22 PEArray.scala 60:13]
  wire [15:0] _GEN_7 = 6'h1 == L0Index ? L0Memory_1 : L0Memory_0; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_8 = 6'h2 == L0Index ? L0Memory_2 : _GEN_7; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_9 = 6'h3 == L0Index ? L0Memory_3 : _GEN_8; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_10 = 6'h4 == L0Index ? L0Memory_4 : _GEN_9; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_11 = 6'h5 == L0Index ? L0Memory_5 : _GEN_10; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_12 = 6'h6 == L0Index ? L0Memory_6 : _GEN_11; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_13 = 6'h7 == L0Index ? L0Memory_7 : _GEN_12; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_14 = 6'h8 == L0Index ? L0Memory_8 : _GEN_13; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_15 = 6'h9 == L0Index ? L0Memory_9 : _GEN_14; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_16 = 6'ha == L0Index ? L0Memory_10 : _GEN_15; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_17 = 6'hb == L0Index ? L0Memory_11 : _GEN_16; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_18 = 6'hc == L0Index ? L0Memory_12 : _GEN_17; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_19 = 6'hd == L0Index ? L0Memory_13 : _GEN_18; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_20 = 6'he == L0Index ? L0Memory_14 : _GEN_19; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_21 = 6'hf == L0Index ? L0Memory_15 : _GEN_20; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_22 = 6'h10 == L0Index ? L0Memory_16 : _GEN_21; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_23 = 6'h11 == L0Index ? L0Memory_17 : _GEN_22; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_24 = 6'h12 == L0Index ? L0Memory_18 : _GEN_23; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_25 = 6'h13 == L0Index ? L0Memory_19 : _GEN_24; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_26 = 6'h14 == L0Index ? L0Memory_20 : _GEN_25; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_27 = 6'h15 == L0Index ? L0Memory_21 : _GEN_26; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_28 = 6'h16 == L0Index ? L0Memory_22 : _GEN_27; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_29 = 6'h17 == L0Index ? L0Memory_23 : _GEN_28; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_30 = 6'h18 == L0Index ? L0Memory_24 : _GEN_29; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_31 = 6'h19 == L0Index ? L0Memory_25 : _GEN_30; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_32 = 6'h1a == L0Index ? L0Memory_26 : _GEN_31; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_33 = 6'h1b == L0Index ? L0Memory_27 : _GEN_32; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_34 = 6'h1c == L0Index ? L0Memory_28 : _GEN_33; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_35 = 6'h1d == L0Index ? L0Memory_29 : _GEN_34; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_36 = 6'h1e == L0Index ? L0Memory_30 : _GEN_35; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_37 = 6'h1f == L0Index ? L0Memory_31 : _GEN_36; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_38 = 6'h20 == L0Index ? L0Memory_32 : _GEN_37; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_39 = 6'h21 == L0Index ? L0Memory_33 : _GEN_38; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_40 = 6'h22 == L0Index ? L0Memory_34 : _GEN_39; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_41 = 6'h23 == L0Index ? L0Memory_35 : _GEN_40; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_42 = 6'h24 == L0Index ? L0Memory_36 : _GEN_41; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_43 = 6'h25 == L0Index ? L0Memory_37 : _GEN_42; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_44 = 6'h26 == L0Index ? L0Memory_38 : _GEN_43; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_45 = 6'h27 == L0Index ? L0Memory_39 : _GEN_44; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_46 = 6'h28 == L0Index ? L0Memory_40 : _GEN_45; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_47 = 6'h29 == L0Index ? L0Memory_41 : _GEN_46; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_48 = 6'h2a == L0Index ? L0Memory_42 : _GEN_47; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_49 = 6'h2b == L0Index ? L0Memory_43 : _GEN_48; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_50 = 6'h2c == L0Index ? L0Memory_44 : _GEN_49; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_51 = 6'h2d == L0Index ? L0Memory_45 : _GEN_50; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_52 = 6'h2e == L0Index ? L0Memory_46 : _GEN_51; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_53 = 6'h2f == L0Index ? L0Memory_47 : _GEN_52; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_54 = 6'h30 == L0Index ? L0Memory_48 : _GEN_53; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_55 = 6'h31 == L0Index ? L0Memory_49 : _GEN_54; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_56 = 6'h32 == L0Index ? L0Memory_50 : _GEN_55; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_57 = 6'h33 == L0Index ? L0Memory_51 : _GEN_56; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_58 = 6'h34 == L0Index ? L0Memory_52 : _GEN_57; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_59 = 6'h35 == L0Index ? L0Memory_53 : _GEN_58; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_60 = 6'h36 == L0Index ? L0Memory_54 : _GEN_59; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_61 = 6'h37 == L0Index ? L0Memory_55 : _GEN_60; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_62 = 6'h38 == L0Index ? L0Memory_56 : _GEN_61; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_63 = 6'h39 == L0Index ? L0Memory_57 : _GEN_62; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_64 = 6'h3a == L0Index ? L0Memory_58 : _GEN_63; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_65 = 6'h3b == L0Index ? L0Memory_59 : _GEN_64; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_66 = 6'h3c == L0Index ? L0Memory_60 : _GEN_65; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_67 = 6'h3d == L0Index ? L0Memory_61 : _GEN_66; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_68 = 6'h3e == L0Index ? L0Memory_62 : _GEN_67; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_69 = 6'h3f == L0Index ? L0Memory_63 : _GEN_68; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [6:0] _GEN_793 = {{1'd0}, L0Index}; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_70 = 7'h40 == _GEN_793 ? L0Memory_64 : _GEN_69; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_71 = 7'h41 == _GEN_793 ? L0Memory_65 : _GEN_70; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_72 = 7'h42 == _GEN_793 ? L0Memory_66 : _GEN_71; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_73 = 7'h43 == _GEN_793 ? L0Memory_67 : _GEN_72; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_74 = 7'h44 == _GEN_793 ? L0Memory_68 : _GEN_73; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_75 = 7'h45 == _GEN_793 ? L0Memory_69 : _GEN_74; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_76 = 7'h46 == _GEN_793 ? L0Memory_70 : _GEN_75; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_77 = 7'h47 == _GEN_793 ? L0Memory_71 : _GEN_76; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_78 = 7'h48 == _GEN_793 ? L0Memory_72 : _GEN_77; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_79 = 7'h49 == _GEN_793 ? L0Memory_73 : _GEN_78; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_80 = 7'h4a == _GEN_793 ? L0Memory_74 : _GEN_79; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_81 = 7'h4b == _GEN_793 ? L0Memory_75 : _GEN_80; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_82 = 7'h4c == _GEN_793 ? L0Memory_76 : _GEN_81; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_83 = 7'h4d == _GEN_793 ? L0Memory_77 : _GEN_82; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_84 = 7'h4e == _GEN_793 ? L0Memory_78 : _GEN_83; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_85 = 7'h4f == _GEN_793 ? L0Memory_79 : _GEN_84; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_86 = 7'h50 == _GEN_793 ? L0Memory_80 : _GEN_85; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_87 = 7'h51 == _GEN_793 ? L0Memory_81 : _GEN_86; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_88 = 7'h52 == _GEN_793 ? L0Memory_82 : _GEN_87; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_89 = 7'h53 == _GEN_793 ? L0Memory_83 : _GEN_88; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_90 = 7'h54 == _GEN_793 ? L0Memory_84 : _GEN_89; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_91 = 7'h55 == _GEN_793 ? L0Memory_85 : _GEN_90; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_92 = 7'h56 == _GEN_793 ? L0Memory_86 : _GEN_91; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_93 = 7'h57 == _GEN_793 ? L0Memory_87 : _GEN_92; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_94 = 7'h58 == _GEN_793 ? L0Memory_88 : _GEN_93; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_95 = 7'h59 == _GEN_793 ? L0Memory_89 : _GEN_94; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_96 = 7'h5a == _GEN_793 ? L0Memory_90 : _GEN_95; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_97 = 7'h5b == _GEN_793 ? L0Memory_91 : _GEN_96; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_98 = 7'h5c == _GEN_793 ? L0Memory_92 : _GEN_97; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_99 = 7'h5d == _GEN_793 ? L0Memory_93 : _GEN_98; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_100 = 7'h5e == _GEN_793 ? L0Memory_94 : _GEN_99; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_101 = 7'h5f == _GEN_793 ? L0Memory_95 : _GEN_100; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_102 = 7'h60 == _GEN_793 ? L0Memory_96 : _GEN_101; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_103 = 7'h61 == _GEN_793 ? L0Memory_97 : _GEN_102; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_104 = 7'h62 == _GEN_793 ? L0Memory_98 : _GEN_103; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_105 = 7'h63 == _GEN_793 ? L0Memory_99 : _GEN_104; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire  _GEN_575 = _T_12 ? 1'h0 : _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 157:12]
  wire  sel5 = _T_3 ? 1'h0 : _GEN_575; // @[Conditional.scala 40:58 PEArray.scala 112:12]
  reg [15:0] mux2out_reg; // @[PEArray.scala 90:28]
  reg [15:0] mux3out_reg; // @[PEArray.scala 91:28]
  reg [9:0] count; // @[PEArray.scala 101:22]
  reg [5:0] GRU_out_width; // @[PEArray.scala 104:26]
  wire [7:0] _GEN_118 = io_control_signal_mask[1] ? 8'h0 : {{2'd0}, GRU_out_width}; // @[PEArray.scala 116:57 PEArray.scala 145:23 PEArray.scala 104:26]
  wire [9:0] _count_T_1 = count + 10'h1; // @[PEArray.scala 162:24]
  wire [9:0] _GEN_120 = count != 10'h33 ? _count_T_1 : count; // @[PEArray.scala 161:27 PEArray.scala 162:15 PEArray.scala 101:22]
  wire [9:0] _GEN_124 = count != 10'h188 ? _count_T_1 : count; // @[PEArray.scala 183:28 PEArray.scala 184:15 PEArray.scala 101:22]
  wire [9:0] _GEN_125 = count == 10'h188 ? 10'h0 : _GEN_124; // @[PEArray.scala 186:28 PEArray.scala 187:15]
  wire [2:0] _GEN_126 = count == 10'h188 ? 3'h0 : state; // @[PEArray.scala 186:28 PEArray.scala 188:15 PEArray.scala 100:22]
  wire [9:0] _GEN_127 = count != 10'h0 ? _count_T_1 : count; // @[PEArray.scala 192:32 PEArray.scala 193:15 PEArray.scala 101:22]
  wire  _T_24 = count == 10'h0; // @[PEArray.scala 195:18]
  wire [5:0] _GEN_128 = count == 10'h0 ? 6'h0 : L0Index; // @[PEArray.scala 195:26 PEArray.scala 196:17 PEArray.scala 39:24]
  wire [9:0] _T_27 = 10'h0 - 10'h1; // @[PEArray.scala 198:51]
  wire [15:0] _GEN_129 = 6'h0 == L0Index ? io_FromL1 : L0Memory_0; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_130 = 6'h1 == L0Index ? io_FromL1 : L0Memory_1; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_131 = 6'h2 == L0Index ? io_FromL1 : L0Memory_2; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_132 = 6'h3 == L0Index ? io_FromL1 : L0Memory_3; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_133 = 6'h4 == L0Index ? io_FromL1 : L0Memory_4; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_134 = 6'h5 == L0Index ? io_FromL1 : L0Memory_5; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_135 = 6'h6 == L0Index ? io_FromL1 : L0Memory_6; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_136 = 6'h7 == L0Index ? io_FromL1 : L0Memory_7; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_137 = 6'h8 == L0Index ? io_FromL1 : L0Memory_8; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_138 = 6'h9 == L0Index ? io_FromL1 : L0Memory_9; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_139 = 6'ha == L0Index ? io_FromL1 : L0Memory_10; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_140 = 6'hb == L0Index ? io_FromL1 : L0Memory_11; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_141 = 6'hc == L0Index ? io_FromL1 : L0Memory_12; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_142 = 6'hd == L0Index ? io_FromL1 : L0Memory_13; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_143 = 6'he == L0Index ? io_FromL1 : L0Memory_14; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_144 = 6'hf == L0Index ? io_FromL1 : L0Memory_15; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_145 = 6'h10 == L0Index ? io_FromL1 : L0Memory_16; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_146 = 6'h11 == L0Index ? io_FromL1 : L0Memory_17; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_147 = 6'h12 == L0Index ? io_FromL1 : L0Memory_18; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_148 = 6'h13 == L0Index ? io_FromL1 : L0Memory_19; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_149 = 6'h14 == L0Index ? io_FromL1 : L0Memory_20; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_150 = 6'h15 == L0Index ? io_FromL1 : L0Memory_21; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_151 = 6'h16 == L0Index ? io_FromL1 : L0Memory_22; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_152 = 6'h17 == L0Index ? io_FromL1 : L0Memory_23; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_153 = 6'h18 == L0Index ? io_FromL1 : L0Memory_24; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_154 = 6'h19 == L0Index ? io_FromL1 : L0Memory_25; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_155 = 6'h1a == L0Index ? io_FromL1 : L0Memory_26; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_156 = 6'h1b == L0Index ? io_FromL1 : L0Memory_27; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_157 = 6'h1c == L0Index ? io_FromL1 : L0Memory_28; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_158 = 6'h1d == L0Index ? io_FromL1 : L0Memory_29; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_159 = 6'h1e == L0Index ? io_FromL1 : L0Memory_30; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_160 = 6'h1f == L0Index ? io_FromL1 : L0Memory_31; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_161 = 6'h20 == L0Index ? io_FromL1 : L0Memory_32; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_162 = 6'h21 == L0Index ? io_FromL1 : L0Memory_33; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_163 = 6'h22 == L0Index ? io_FromL1 : L0Memory_34; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_164 = 6'h23 == L0Index ? io_FromL1 : L0Memory_35; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_165 = 6'h24 == L0Index ? io_FromL1 : L0Memory_36; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_166 = 6'h25 == L0Index ? io_FromL1 : L0Memory_37; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_167 = 6'h26 == L0Index ? io_FromL1 : L0Memory_38; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_168 = 6'h27 == L0Index ? io_FromL1 : L0Memory_39; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_169 = 6'h28 == L0Index ? io_FromL1 : L0Memory_40; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_170 = 6'h29 == L0Index ? io_FromL1 : L0Memory_41; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_171 = 6'h2a == L0Index ? io_FromL1 : L0Memory_42; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_172 = 6'h2b == L0Index ? io_FromL1 : L0Memory_43; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_173 = 6'h2c == L0Index ? io_FromL1 : L0Memory_44; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_174 = 6'h2d == L0Index ? io_FromL1 : L0Memory_45; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_175 = 6'h2e == L0Index ? io_FromL1 : L0Memory_46; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_176 = 6'h2f == L0Index ? io_FromL1 : L0Memory_47; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_177 = 6'h30 == L0Index ? io_FromL1 : L0Memory_48; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_178 = 6'h31 == L0Index ? io_FromL1 : L0Memory_49; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_179 = 6'h32 == L0Index ? io_FromL1 : L0Memory_50; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_180 = 6'h33 == L0Index ? io_FromL1 : L0Memory_51; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_181 = 6'h34 == L0Index ? io_FromL1 : L0Memory_52; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_182 = 6'h35 == L0Index ? io_FromL1 : L0Memory_53; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_183 = 6'h36 == L0Index ? io_FromL1 : L0Memory_54; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_184 = 6'h37 == L0Index ? io_FromL1 : L0Memory_55; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_185 = 6'h38 == L0Index ? io_FromL1 : L0Memory_56; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_186 = 6'h39 == L0Index ? io_FromL1 : L0Memory_57; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_187 = 6'h3a == L0Index ? io_FromL1 : L0Memory_58; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_188 = 6'h3b == L0Index ? io_FromL1 : L0Memory_59; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_189 = 6'h3c == L0Index ? io_FromL1 : L0Memory_60; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_190 = 6'h3d == L0Index ? io_FromL1 : L0Memory_61; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_191 = 6'h3e == L0Index ? io_FromL1 : L0Memory_62; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_192 = 6'h3f == L0Index ? io_FromL1 : L0Memory_63; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_193 = 7'h40 == _GEN_793 ? io_FromL1 : L0Memory_64; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_194 = 7'h41 == _GEN_793 ? io_FromL1 : L0Memory_65; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_195 = 7'h42 == _GEN_793 ? io_FromL1 : L0Memory_66; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_196 = 7'h43 == _GEN_793 ? io_FromL1 : L0Memory_67; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_197 = 7'h44 == _GEN_793 ? io_FromL1 : L0Memory_68; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_198 = 7'h45 == _GEN_793 ? io_FromL1 : L0Memory_69; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_199 = 7'h46 == _GEN_793 ? io_FromL1 : L0Memory_70; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_200 = 7'h47 == _GEN_793 ? io_FromL1 : L0Memory_71; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_201 = 7'h48 == _GEN_793 ? io_FromL1 : L0Memory_72; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_202 = 7'h49 == _GEN_793 ? io_FromL1 : L0Memory_73; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_203 = 7'h4a == _GEN_793 ? io_FromL1 : L0Memory_74; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_204 = 7'h4b == _GEN_793 ? io_FromL1 : L0Memory_75; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_205 = 7'h4c == _GEN_793 ? io_FromL1 : L0Memory_76; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_206 = 7'h4d == _GEN_793 ? io_FromL1 : L0Memory_77; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_207 = 7'h4e == _GEN_793 ? io_FromL1 : L0Memory_78; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_208 = 7'h4f == _GEN_793 ? io_FromL1 : L0Memory_79; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_209 = 7'h50 == _GEN_793 ? io_FromL1 : L0Memory_80; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_210 = 7'h51 == _GEN_793 ? io_FromL1 : L0Memory_81; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_211 = 7'h52 == _GEN_793 ? io_FromL1 : L0Memory_82; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_212 = 7'h53 == _GEN_793 ? io_FromL1 : L0Memory_83; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_213 = 7'h54 == _GEN_793 ? io_FromL1 : L0Memory_84; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_214 = 7'h55 == _GEN_793 ? io_FromL1 : L0Memory_85; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_215 = 7'h56 == _GEN_793 ? io_FromL1 : L0Memory_86; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_216 = 7'h57 == _GEN_793 ? io_FromL1 : L0Memory_87; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_217 = 7'h58 == _GEN_793 ? io_FromL1 : L0Memory_88; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_218 = 7'h59 == _GEN_793 ? io_FromL1 : L0Memory_89; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_219 = 7'h5a == _GEN_793 ? io_FromL1 : L0Memory_90; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_220 = 7'h5b == _GEN_793 ? io_FromL1 : L0Memory_91; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_221 = 7'h5c == _GEN_793 ? io_FromL1 : L0Memory_92; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_222 = 7'h5d == _GEN_793 ? io_FromL1 : L0Memory_93; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_223 = 7'h5e == _GEN_793 ? io_FromL1 : L0Memory_94; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_224 = 7'h5f == _GEN_793 ? io_FromL1 : L0Memory_95; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_225 = 7'h60 == _GEN_793 ? io_FromL1 : L0Memory_96; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_226 = 7'h61 == _GEN_793 ? io_FromL1 : L0Memory_97; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_227 = 7'h62 == _GEN_793 ? io_FromL1 : L0Memory_98; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_228 = 7'h63 == _GEN_793 ? io_FromL1 : L0Memory_99; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [5:0] _L0Index_T_2 = L0Index + 6'h1; // @[PEArray.scala 200:28]
  wire [15:0] _GEN_229 = count >= 10'h1 & count <= _T_27 ? _GEN_129 : L0Memory_0; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_230 = count >= 10'h1 & count <= _T_27 ? _GEN_130 : L0Memory_1; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_231 = count >= 10'h1 & count <= _T_27 ? _GEN_131 : L0Memory_2; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_232 = count >= 10'h1 & count <= _T_27 ? _GEN_132 : L0Memory_3; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_233 = count >= 10'h1 & count <= _T_27 ? _GEN_133 : L0Memory_4; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_234 = count >= 10'h1 & count <= _T_27 ? _GEN_134 : L0Memory_5; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_235 = count >= 10'h1 & count <= _T_27 ? _GEN_135 : L0Memory_6; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_236 = count >= 10'h1 & count <= _T_27 ? _GEN_136 : L0Memory_7; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_237 = count >= 10'h1 & count <= _T_27 ? _GEN_137 : L0Memory_8; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_238 = count >= 10'h1 & count <= _T_27 ? _GEN_138 : L0Memory_9; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_239 = count >= 10'h1 & count <= _T_27 ? _GEN_139 : L0Memory_10; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_240 = count >= 10'h1 & count <= _T_27 ? _GEN_140 : L0Memory_11; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_241 = count >= 10'h1 & count <= _T_27 ? _GEN_141 : L0Memory_12; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_242 = count >= 10'h1 & count <= _T_27 ? _GEN_142 : L0Memory_13; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_243 = count >= 10'h1 & count <= _T_27 ? _GEN_143 : L0Memory_14; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_244 = count >= 10'h1 & count <= _T_27 ? _GEN_144 : L0Memory_15; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_245 = count >= 10'h1 & count <= _T_27 ? _GEN_145 : L0Memory_16; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_246 = count >= 10'h1 & count <= _T_27 ? _GEN_146 : L0Memory_17; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_247 = count >= 10'h1 & count <= _T_27 ? _GEN_147 : L0Memory_18; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_248 = count >= 10'h1 & count <= _T_27 ? _GEN_148 : L0Memory_19; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_249 = count >= 10'h1 & count <= _T_27 ? _GEN_149 : L0Memory_20; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_250 = count >= 10'h1 & count <= _T_27 ? _GEN_150 : L0Memory_21; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_251 = count >= 10'h1 & count <= _T_27 ? _GEN_151 : L0Memory_22; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_252 = count >= 10'h1 & count <= _T_27 ? _GEN_152 : L0Memory_23; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_253 = count >= 10'h1 & count <= _T_27 ? _GEN_153 : L0Memory_24; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_254 = count >= 10'h1 & count <= _T_27 ? _GEN_154 : L0Memory_25; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_255 = count >= 10'h1 & count <= _T_27 ? _GEN_155 : L0Memory_26; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_256 = count >= 10'h1 & count <= _T_27 ? _GEN_156 : L0Memory_27; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_257 = count >= 10'h1 & count <= _T_27 ? _GEN_157 : L0Memory_28; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_258 = count >= 10'h1 & count <= _T_27 ? _GEN_158 : L0Memory_29; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_259 = count >= 10'h1 & count <= _T_27 ? _GEN_159 : L0Memory_30; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_260 = count >= 10'h1 & count <= _T_27 ? _GEN_160 : L0Memory_31; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_261 = count >= 10'h1 & count <= _T_27 ? _GEN_161 : L0Memory_32; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_262 = count >= 10'h1 & count <= _T_27 ? _GEN_162 : L0Memory_33; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_263 = count >= 10'h1 & count <= _T_27 ? _GEN_163 : L0Memory_34; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_264 = count >= 10'h1 & count <= _T_27 ? _GEN_164 : L0Memory_35; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_265 = count >= 10'h1 & count <= _T_27 ? _GEN_165 : L0Memory_36; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_266 = count >= 10'h1 & count <= _T_27 ? _GEN_166 : L0Memory_37; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_267 = count >= 10'h1 & count <= _T_27 ? _GEN_167 : L0Memory_38; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_268 = count >= 10'h1 & count <= _T_27 ? _GEN_168 : L0Memory_39; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_269 = count >= 10'h1 & count <= _T_27 ? _GEN_169 : L0Memory_40; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_270 = count >= 10'h1 & count <= _T_27 ? _GEN_170 : L0Memory_41; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_271 = count >= 10'h1 & count <= _T_27 ? _GEN_171 : L0Memory_42; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_272 = count >= 10'h1 & count <= _T_27 ? _GEN_172 : L0Memory_43; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_273 = count >= 10'h1 & count <= _T_27 ? _GEN_173 : L0Memory_44; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_274 = count >= 10'h1 & count <= _T_27 ? _GEN_174 : L0Memory_45; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_275 = count >= 10'h1 & count <= _T_27 ? _GEN_175 : L0Memory_46; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_276 = count >= 10'h1 & count <= _T_27 ? _GEN_176 : L0Memory_47; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_277 = count >= 10'h1 & count <= _T_27 ? _GEN_177 : L0Memory_48; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_278 = count >= 10'h1 & count <= _T_27 ? _GEN_178 : L0Memory_49; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_279 = count >= 10'h1 & count <= _T_27 ? _GEN_179 : L0Memory_50; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_280 = count >= 10'h1 & count <= _T_27 ? _GEN_180 : L0Memory_51; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_281 = count >= 10'h1 & count <= _T_27 ? _GEN_181 : L0Memory_52; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_282 = count >= 10'h1 & count <= _T_27 ? _GEN_182 : L0Memory_53; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_283 = count >= 10'h1 & count <= _T_27 ? _GEN_183 : L0Memory_54; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_284 = count >= 10'h1 & count <= _T_27 ? _GEN_184 : L0Memory_55; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_285 = count >= 10'h1 & count <= _T_27 ? _GEN_185 : L0Memory_56; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_286 = count >= 10'h1 & count <= _T_27 ? _GEN_186 : L0Memory_57; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_287 = count >= 10'h1 & count <= _T_27 ? _GEN_187 : L0Memory_58; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_288 = count >= 10'h1 & count <= _T_27 ? _GEN_188 : L0Memory_59; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_289 = count >= 10'h1 & count <= _T_27 ? _GEN_189 : L0Memory_60; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_290 = count >= 10'h1 & count <= _T_27 ? _GEN_190 : L0Memory_61; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_291 = count >= 10'h1 & count <= _T_27 ? _GEN_191 : L0Memory_62; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_292 = count >= 10'h1 & count <= _T_27 ? _GEN_192 : L0Memory_63; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_293 = count >= 10'h1 & count <= _T_27 ? _GEN_193 : L0Memory_64; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_294 = count >= 10'h1 & count <= _T_27 ? _GEN_194 : L0Memory_65; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_295 = count >= 10'h1 & count <= _T_27 ? _GEN_195 : L0Memory_66; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_296 = count >= 10'h1 & count <= _T_27 ? _GEN_196 : L0Memory_67; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_297 = count >= 10'h1 & count <= _T_27 ? _GEN_197 : L0Memory_68; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_298 = count >= 10'h1 & count <= _T_27 ? _GEN_198 : L0Memory_69; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_299 = count >= 10'h1 & count <= _T_27 ? _GEN_199 : L0Memory_70; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_300 = count >= 10'h1 & count <= _T_27 ? _GEN_200 : L0Memory_71; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_301 = count >= 10'h1 & count <= _T_27 ? _GEN_201 : L0Memory_72; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_302 = count >= 10'h1 & count <= _T_27 ? _GEN_202 : L0Memory_73; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_303 = count >= 10'h1 & count <= _T_27 ? _GEN_203 : L0Memory_74; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_304 = count >= 10'h1 & count <= _T_27 ? _GEN_204 : L0Memory_75; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_305 = count >= 10'h1 & count <= _T_27 ? _GEN_205 : L0Memory_76; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_306 = count >= 10'h1 & count <= _T_27 ? _GEN_206 : L0Memory_77; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_307 = count >= 10'h1 & count <= _T_27 ? _GEN_207 : L0Memory_78; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_308 = count >= 10'h1 & count <= _T_27 ? _GEN_208 : L0Memory_79; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_309 = count >= 10'h1 & count <= _T_27 ? _GEN_209 : L0Memory_80; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_310 = count >= 10'h1 & count <= _T_27 ? _GEN_210 : L0Memory_81; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_311 = count >= 10'h1 & count <= _T_27 ? _GEN_211 : L0Memory_82; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_312 = count >= 10'h1 & count <= _T_27 ? _GEN_212 : L0Memory_83; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_313 = count >= 10'h1 & count <= _T_27 ? _GEN_213 : L0Memory_84; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_314 = count >= 10'h1 & count <= _T_27 ? _GEN_214 : L0Memory_85; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_315 = count >= 10'h1 & count <= _T_27 ? _GEN_215 : L0Memory_86; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_316 = count >= 10'h1 & count <= _T_27 ? _GEN_216 : L0Memory_87; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_317 = count >= 10'h1 & count <= _T_27 ? _GEN_217 : L0Memory_88; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_318 = count >= 10'h1 & count <= _T_27 ? _GEN_218 : L0Memory_89; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_319 = count >= 10'h1 & count <= _T_27 ? _GEN_219 : L0Memory_90; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_320 = count >= 10'h1 & count <= _T_27 ? _GEN_220 : L0Memory_91; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_321 = count >= 10'h1 & count <= _T_27 ? _GEN_221 : L0Memory_92; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_322 = count >= 10'h1 & count <= _T_27 ? _GEN_222 : L0Memory_93; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_323 = count >= 10'h1 & count <= _T_27 ? _GEN_223 : L0Memory_94; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_324 = count >= 10'h1 & count <= _T_27 ? _GEN_224 : L0Memory_95; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_325 = count >= 10'h1 & count <= _T_27 ? _GEN_225 : L0Memory_96; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_326 = count >= 10'h1 & count <= _T_27 ? _GEN_226 : L0Memory_97; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_327 = count >= 10'h1 & count <= _T_27 ? _GEN_227 : L0Memory_98; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_328 = count >= 10'h1 & count <= _T_27 ? _GEN_228 : L0Memory_99; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [5:0] _GEN_329 = count >= 10'h1 & count <= _T_27 ? _L0Index_T_2 : _GEN_128; // @[PEArray.scala 198:59 PEArray.scala 200:17]
  wire [9:0] _GEN_330 = _T_24 ? 10'h0 : _GEN_127; // @[PEArray.scala 202:32 PEArray.scala 203:15]
  wire [2:0] _GEN_331 = _T_24 ? 3'h0 : state; // @[PEArray.scala 202:32 PEArray.scala 204:15 PEArray.scala 100:22]
  wire [9:0] _GEN_865 = {{4'd0}, GRU_out_width}; // @[PEArray.scala 220:19]
  wire [9:0] _GEN_0 = count % _GEN_865; // @[PEArray.scala 220:19]
  wire [5:0] _T_36 = _GEN_0[5:0]; // @[PEArray.scala 220:19]
  wire [5:0] _T_38 = GRU_out_width - 6'h1; // @[PEArray.scala 220:55]
  wire [5:0] _GEN_334 = _T_36 == _T_38 ? _L0Index_T_2 : 6'h0; // @[PEArray.scala 220:62 PEArray.scala 221:17 PEArray.scala 214:15]
  wire [5:0] _GEN_346 = _T_41 ? _GEN_334 : L0Index; // @[Conditional.scala 39:67 PEArray.scala 39:24]
  wire [9:0] _GEN_347 = _T_41 ? _GEN_330 : count; // @[Conditional.scala 39:67 PEArray.scala 101:22]
  wire [2:0] _GEN_348 = _T_41 ? _GEN_331 : state; // @[Conditional.scala 39:67 PEArray.scala 100:22]
  wire [5:0] _GEN_353 = _T_31 ? _GEN_334 : _GEN_346; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_354 = _T_31 ? _GEN_330 : _GEN_347; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_355 = _T_31 ? _GEN_331 : _GEN_348; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_356 = _T_22 ? _GEN_330 : _GEN_354; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_357 = _T_22 ? _GEN_329 : _GEN_353; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_458 = _T_22 ? _GEN_331 : _GEN_355; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_690 = _T_3 ? _GEN_118 : {{2'd0}, GRU_out_width}; // @[Conditional.scala 40:58 PEArray.scala 104:26]
  FP16MulAdder FP16MAC ( // @[PEArray.scala 72:23]
    .io_a(FP16MAC_io_a),
    .io_b(FP16MAC_io_b),
    .io_c(FP16MAC_io_c),
    .io_out(FP16MAC_io_out)
  );
  assign io_ToRightPE = mux3out_reg; // @[PEArray.scala 95:16]
  assign io_ToBelowPE = mux2out_reg; // @[PEArray.scala 94:16]
  assign FP16MAC_io_a = sel1 ? io_FromL1 : io_FromLeftPE; // @[PEArray.scala 50:14 PEArray.scala 50:23 PEArray.scala 51:24]
  assign FP16MAC_io_b = sel5 ? mux4out : _GEN_105; // @[PEArray.scala 77:13 PEArray.scala 78:18 PEArray.scala 81:18]
  assign FP16MAC_io_c = sel5 ? _GEN_105 : mux4out; // @[PEArray.scala 77:13 PEArray.scala 79:18 PEArray.scala 82:18]
  always @(posedge clock) begin
    if (reset) begin // @[PEArray.scala 39:24]
      L0Index <= 6'h0; // @[PEArray.scala 39:24]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h0; // @[PEArray.scala 159:15]
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        L0Index <= 6'hd; // @[PEArray.scala 181:15]
      end else begin
        L0Index <= _GEN_357;
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_0 <= _GEN_229;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_1 <= _GEN_230;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_2 <= _GEN_231;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_3 <= _GEN_232;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_4 <= _GEN_233;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_5 <= _GEN_234;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_6 <= _GEN_235;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_7 <= _GEN_236;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_8 <= _GEN_237;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_9 <= _GEN_238;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_10 <= _GEN_239;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_11 <= _GEN_240;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_12 <= _GEN_241;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_13 <= _GEN_242;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_14 <= _GEN_243;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_15 <= _GEN_244;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_16 <= _GEN_245;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_17 <= _GEN_246;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_18 <= _GEN_247;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_19 <= _GEN_248;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_20 <= _GEN_249;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_21 <= _GEN_250;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_22 <= _GEN_251;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_23 <= _GEN_252;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_24 <= _GEN_253;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_25 <= _GEN_254;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_26 <= _GEN_255;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_27 <= _GEN_256;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_28 <= _GEN_257;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_29 <= _GEN_258;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_30 <= _GEN_259;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_31 <= _GEN_260;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_32 <= _GEN_261;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_33 <= _GEN_262;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_34 <= _GEN_263;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_35 <= _GEN_264;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_36 <= _GEN_265;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_37 <= _GEN_266;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_38 <= _GEN_267;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_39 <= _GEN_268;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_40 <= _GEN_269;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_41 <= _GEN_270;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_42 <= _GEN_271;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_43 <= _GEN_272;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_44 <= _GEN_273;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_45 <= _GEN_274;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_46 <= _GEN_275;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_47 <= _GEN_276;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_48 <= _GEN_277;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_49 <= _GEN_278;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_50 <= _GEN_279;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_51 <= _GEN_280;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_52 <= _GEN_281;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_53 <= _GEN_282;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_54 <= _GEN_283;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_55 <= _GEN_284;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_56 <= _GEN_285;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_57 <= _GEN_286;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_58 <= _GEN_287;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_59 <= _GEN_288;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_60 <= _GEN_289;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_61 <= _GEN_290;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_62 <= _GEN_291;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_63 <= _GEN_292;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_64 <= _GEN_293;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_65 <= _GEN_294;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_66 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_67 <= _GEN_296;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_68 <= _GEN_297;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_69 <= _GEN_298;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_70 <= _GEN_299;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_71 <= _GEN_300;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_72 <= _GEN_301;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_73 <= _GEN_302;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_74 <= _GEN_303;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_75 <= _GEN_304;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_76 <= _GEN_305;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_77 <= _GEN_306;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_78 <= _GEN_307;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_79 <= _GEN_308;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_80 <= _GEN_309;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_81 <= _GEN_310;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_82 <= _GEN_311;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_83 <= _GEN_312;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_84 <= _GEN_313;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_85 <= _GEN_314;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_86 <= _GEN_315;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_87 <= _GEN_316;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_88 <= _GEN_317;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_89 <= _GEN_318;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_90 <= _GEN_319;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_91 <= _GEN_320;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_92 <= _GEN_321;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_93 <= _GEN_322;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_94 <= _GEN_323;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_95 <= _GEN_324;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_96 <= _GEN_325;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_97 <= _GEN_326;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_98 <= _GEN_327;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_99 <= _GEN_328;
          end
        end
      end
    end
    if (reset) begin // @[PEArray.scala 100:22]
      state <= 3'h0; // @[PEArray.scala 100:22]
    end else if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[1]) begin // @[PEArray.scala 116:57]
        state <= 3'h1;
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      if (count == 10'h33) begin // @[PEArray.scala 164:27]
        state <= 3'h0; // @[PEArray.scala 166:15]
      end
    end else if (_T_16) begin // @[Conditional.scala 39:67]
      state <= _GEN_126;
    end else begin
      state <= _GEN_458;
    end
    if (reset) begin // @[PEArray.scala 90:28]
      mux2out_reg <= 16'h0; // @[PEArray.scala 90:28]
    end else begin
      mux2out_reg <= MAC_out; // @[PEArray.scala 90:28]
    end
    if (reset) begin // @[PEArray.scala 91:28]
      mux3out_reg <= 16'h0; // @[PEArray.scala 91:28]
    end else if (sel3) begin // @[PEArray.scala 56:14]
      mux3out_reg <= MAC_out; // @[PEArray.scala 56:23]
    end else if (sel1) begin // @[PEArray.scala 50:14]
      mux3out_reg <= io_FromL1; // @[PEArray.scala 50:23]
    end else begin
      mux3out_reg <= io_FromLeftPE; // @[PEArray.scala 51:24]
    end
    if (reset) begin // @[PEArray.scala 101:22]
      count <= 10'h0; // @[PEArray.scala 101:22]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        if (count == 10'h33) begin // @[PEArray.scala 164:27]
          count <= 10'h0; // @[PEArray.scala 165:15]
        end else begin
          count <= _GEN_120;
        end
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        count <= _GEN_125;
      end else begin
        count <= _GEN_356;
      end
    end
    GRU_out_width <= _GEN_690[5:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  L0Index = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  L0Memory_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  L0Memory_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  L0Memory_2 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  L0Memory_3 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  L0Memory_4 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  L0Memory_5 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  L0Memory_6 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  L0Memory_7 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  L0Memory_8 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  L0Memory_9 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  L0Memory_10 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  L0Memory_11 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  L0Memory_12 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  L0Memory_13 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  L0Memory_14 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  L0Memory_15 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  L0Memory_16 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  L0Memory_17 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  L0Memory_18 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  L0Memory_19 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  L0Memory_20 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  L0Memory_21 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  L0Memory_22 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  L0Memory_23 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  L0Memory_24 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  L0Memory_25 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  L0Memory_26 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  L0Memory_27 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  L0Memory_28 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  L0Memory_29 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  L0Memory_30 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  L0Memory_31 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  L0Memory_32 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  L0Memory_33 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  L0Memory_34 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  L0Memory_35 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  L0Memory_36 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  L0Memory_37 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  L0Memory_38 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  L0Memory_39 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  L0Memory_40 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  L0Memory_41 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  L0Memory_42 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  L0Memory_43 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  L0Memory_44 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  L0Memory_45 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  L0Memory_46 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  L0Memory_47 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  L0Memory_48 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  L0Memory_49 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  L0Memory_50 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  L0Memory_51 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  L0Memory_52 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  L0Memory_53 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  L0Memory_54 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  L0Memory_55 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  L0Memory_56 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  L0Memory_57 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  L0Memory_58 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  L0Memory_59 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  L0Memory_60 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  L0Memory_61 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  L0Memory_62 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  L0Memory_63 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  L0Memory_64 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  L0Memory_65 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  L0Memory_66 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  L0Memory_67 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  L0Memory_68 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  L0Memory_69 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  L0Memory_70 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  L0Memory_71 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  L0Memory_72 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  L0Memory_73 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  L0Memory_74 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  L0Memory_75 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  L0Memory_76 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  L0Memory_77 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  L0Memory_78 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  L0Memory_79 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  L0Memory_80 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  L0Memory_81 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  L0Memory_82 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  L0Memory_83 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  L0Memory_84 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  L0Memory_85 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  L0Memory_86 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  L0Memory_87 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  L0Memory_88 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  L0Memory_89 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  L0Memory_90 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  L0Memory_91 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  L0Memory_92 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  L0Memory_93 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  L0Memory_94 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  L0Memory_95 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  L0Memory_96 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  L0Memory_97 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  L0Memory_98 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  L0Memory_99 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  state = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  mux2out_reg = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  mux3out_reg = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  count = _RAND_104[9:0];
  _RAND_105 = {1{`RANDOM}};
  GRU_out_width = _RAND_105[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PE_31(
  input         clock,
  input         reset,
  input  [15:0] io_FromAbovePE,
  input  [15:0] io_FromLeftPE,
  input  [15:0] io_FromL1,
  input  [11:0] io_control_signal_mask,
  output [15:0] io_ToRightPE,
  output [15:0] io_ToBelowPE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] FP16MAC_io_a; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_b; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_c; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_out; // @[PEArray.scala 72:23]
  reg [5:0] L0Index; // @[PEArray.scala 39:24]
  reg [15:0] L0Memory_0; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_1; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_2; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_3; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_4; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_5; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_6; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_7; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_8; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_9; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_10; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_11; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_12; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_13; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_14; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_15; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_16; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_17; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_18; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_19; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_20; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_21; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_22; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_23; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_24; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_25; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_26; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_27; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_28; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_29; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_30; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_31; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_32; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_33; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_34; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_35; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_36; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_37; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_38; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_39; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_40; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_41; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_42; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_43; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_44; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_45; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_46; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_47; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_48; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_49; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_50; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_51; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_52; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_53; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_54; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_55; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_56; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_57; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_58; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_59; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_60; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_61; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_62; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_63; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_64; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_65; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_66; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_67; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_68; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_69; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_70; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_71; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_72; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_73; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_74; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_75; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_76; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_77; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_78; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_79; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_80; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_81; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_82; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_83; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_84; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_85; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_86; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_87; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_88; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_89; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_90; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_91; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_92; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_93; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_94; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_95; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_96; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_97; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_98; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_99; // @[PEArray.scala 40:21]
  reg [2:0] state; // @[PEArray.scala 100:22]
  wire  _T_3 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_12 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_16 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_22 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_31 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_41 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_342 = _T_41 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 231:12 PEArray.scala 32:8]
  wire  _GEN_349 = _T_31 ? 1'h0 : _GEN_342; // @[Conditional.scala 39:67 PEArray.scala 208:12]
  wire  _GEN_459 = _T_22 | _GEN_349; // @[Conditional.scala 39:67 PEArray.scala 32:8]
  wire  _GEN_463 = _T_16 ? 1'h0 : _GEN_459; // @[Conditional.scala 39:67]
  wire  _GEN_572 = _T_12 | _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 149:12]
  wire  sel1 = _T_3 | _GEN_572; // @[Conditional.scala 40:58 PEArray.scala 108:12]
  wire [15:0] MAC_out = FP16MAC_io_out; // @[PEArray.scala 47:21 PEArray.scala 85:11]
  wire  _GEN_465 = _T_16 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 177:12]
  wire  _GEN_580 = _T_12 | _GEN_465; // @[Conditional.scala 39:67 PEArray.scala 34:8]
  wire  sel3 = _T_3 | _GEN_580; // @[Conditional.scala 40:58 PEArray.scala 110:12]
  wire [1:0] _GEN_344 = _T_41 ? 2'h2 : 2'h0; // @[Conditional.scala 39:67 PEArray.scala 233:12 PEArray.scala 35:8]
  wire [1:0] _GEN_351 = _T_31 ? 2'h2 : _GEN_344; // @[Conditional.scala 39:67 PEArray.scala 210:12]
  wire [1:0] _GEN_461 = _T_22 ? 2'h0 : _GEN_351; // @[Conditional.scala 39:67 PEArray.scala 35:8]
  wire [1:0] _GEN_466 = _T_16 ? 2'h0 : _GEN_461; // @[Conditional.scala 39:67 PEArray.scala 178:12]
  wire [1:0] _GEN_574 = _T_12 ? 2'h1 : _GEN_466; // @[Conditional.scala 39:67]
  wire [1:0] sel4 = _T_3 ? 2'h0 : _GEN_574; // @[Conditional.scala 40:58 PEArray.scala 111:12]
  wire [15:0] _GEN_3 = sel4 == 2'h2 ? io_FromL1 : 16'h0; // @[PEArray.scala 65:28 PEArray.scala 66:15 PEArray.scala 69:15]
  wire [15:0] _GEN_4 = sel4 == 2'h1 ? io_FromAbovePE : _GEN_3; // @[PEArray.scala 62:28 PEArray.scala 63:15]
  wire [15:0] mux4out = sel4 == 2'h0 ? 16'h0 : _GEN_4; // @[PEArray.scala 59:22 PEArray.scala 60:13]
  wire [15:0] _GEN_7 = 6'h1 == L0Index ? L0Memory_1 : L0Memory_0; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_8 = 6'h2 == L0Index ? L0Memory_2 : _GEN_7; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_9 = 6'h3 == L0Index ? L0Memory_3 : _GEN_8; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_10 = 6'h4 == L0Index ? L0Memory_4 : _GEN_9; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_11 = 6'h5 == L0Index ? L0Memory_5 : _GEN_10; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_12 = 6'h6 == L0Index ? L0Memory_6 : _GEN_11; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_13 = 6'h7 == L0Index ? L0Memory_7 : _GEN_12; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_14 = 6'h8 == L0Index ? L0Memory_8 : _GEN_13; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_15 = 6'h9 == L0Index ? L0Memory_9 : _GEN_14; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_16 = 6'ha == L0Index ? L0Memory_10 : _GEN_15; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_17 = 6'hb == L0Index ? L0Memory_11 : _GEN_16; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_18 = 6'hc == L0Index ? L0Memory_12 : _GEN_17; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_19 = 6'hd == L0Index ? L0Memory_13 : _GEN_18; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_20 = 6'he == L0Index ? L0Memory_14 : _GEN_19; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_21 = 6'hf == L0Index ? L0Memory_15 : _GEN_20; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_22 = 6'h10 == L0Index ? L0Memory_16 : _GEN_21; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_23 = 6'h11 == L0Index ? L0Memory_17 : _GEN_22; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_24 = 6'h12 == L0Index ? L0Memory_18 : _GEN_23; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_25 = 6'h13 == L0Index ? L0Memory_19 : _GEN_24; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_26 = 6'h14 == L0Index ? L0Memory_20 : _GEN_25; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_27 = 6'h15 == L0Index ? L0Memory_21 : _GEN_26; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_28 = 6'h16 == L0Index ? L0Memory_22 : _GEN_27; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_29 = 6'h17 == L0Index ? L0Memory_23 : _GEN_28; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_30 = 6'h18 == L0Index ? L0Memory_24 : _GEN_29; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_31 = 6'h19 == L0Index ? L0Memory_25 : _GEN_30; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_32 = 6'h1a == L0Index ? L0Memory_26 : _GEN_31; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_33 = 6'h1b == L0Index ? L0Memory_27 : _GEN_32; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_34 = 6'h1c == L0Index ? L0Memory_28 : _GEN_33; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_35 = 6'h1d == L0Index ? L0Memory_29 : _GEN_34; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_36 = 6'h1e == L0Index ? L0Memory_30 : _GEN_35; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_37 = 6'h1f == L0Index ? L0Memory_31 : _GEN_36; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_38 = 6'h20 == L0Index ? L0Memory_32 : _GEN_37; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_39 = 6'h21 == L0Index ? L0Memory_33 : _GEN_38; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_40 = 6'h22 == L0Index ? L0Memory_34 : _GEN_39; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_41 = 6'h23 == L0Index ? L0Memory_35 : _GEN_40; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_42 = 6'h24 == L0Index ? L0Memory_36 : _GEN_41; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_43 = 6'h25 == L0Index ? L0Memory_37 : _GEN_42; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_44 = 6'h26 == L0Index ? L0Memory_38 : _GEN_43; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_45 = 6'h27 == L0Index ? L0Memory_39 : _GEN_44; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_46 = 6'h28 == L0Index ? L0Memory_40 : _GEN_45; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_47 = 6'h29 == L0Index ? L0Memory_41 : _GEN_46; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_48 = 6'h2a == L0Index ? L0Memory_42 : _GEN_47; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_49 = 6'h2b == L0Index ? L0Memory_43 : _GEN_48; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_50 = 6'h2c == L0Index ? L0Memory_44 : _GEN_49; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_51 = 6'h2d == L0Index ? L0Memory_45 : _GEN_50; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_52 = 6'h2e == L0Index ? L0Memory_46 : _GEN_51; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_53 = 6'h2f == L0Index ? L0Memory_47 : _GEN_52; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_54 = 6'h30 == L0Index ? L0Memory_48 : _GEN_53; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_55 = 6'h31 == L0Index ? L0Memory_49 : _GEN_54; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_56 = 6'h32 == L0Index ? L0Memory_50 : _GEN_55; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_57 = 6'h33 == L0Index ? L0Memory_51 : _GEN_56; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_58 = 6'h34 == L0Index ? L0Memory_52 : _GEN_57; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_59 = 6'h35 == L0Index ? L0Memory_53 : _GEN_58; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_60 = 6'h36 == L0Index ? L0Memory_54 : _GEN_59; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_61 = 6'h37 == L0Index ? L0Memory_55 : _GEN_60; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_62 = 6'h38 == L0Index ? L0Memory_56 : _GEN_61; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_63 = 6'h39 == L0Index ? L0Memory_57 : _GEN_62; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_64 = 6'h3a == L0Index ? L0Memory_58 : _GEN_63; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_65 = 6'h3b == L0Index ? L0Memory_59 : _GEN_64; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_66 = 6'h3c == L0Index ? L0Memory_60 : _GEN_65; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_67 = 6'h3d == L0Index ? L0Memory_61 : _GEN_66; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_68 = 6'h3e == L0Index ? L0Memory_62 : _GEN_67; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_69 = 6'h3f == L0Index ? L0Memory_63 : _GEN_68; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [6:0] _GEN_793 = {{1'd0}, L0Index}; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_70 = 7'h40 == _GEN_793 ? L0Memory_64 : _GEN_69; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_71 = 7'h41 == _GEN_793 ? L0Memory_65 : _GEN_70; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_72 = 7'h42 == _GEN_793 ? L0Memory_66 : _GEN_71; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_73 = 7'h43 == _GEN_793 ? L0Memory_67 : _GEN_72; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_74 = 7'h44 == _GEN_793 ? L0Memory_68 : _GEN_73; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_75 = 7'h45 == _GEN_793 ? L0Memory_69 : _GEN_74; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_76 = 7'h46 == _GEN_793 ? L0Memory_70 : _GEN_75; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_77 = 7'h47 == _GEN_793 ? L0Memory_71 : _GEN_76; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_78 = 7'h48 == _GEN_793 ? L0Memory_72 : _GEN_77; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_79 = 7'h49 == _GEN_793 ? L0Memory_73 : _GEN_78; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_80 = 7'h4a == _GEN_793 ? L0Memory_74 : _GEN_79; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_81 = 7'h4b == _GEN_793 ? L0Memory_75 : _GEN_80; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_82 = 7'h4c == _GEN_793 ? L0Memory_76 : _GEN_81; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_83 = 7'h4d == _GEN_793 ? L0Memory_77 : _GEN_82; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_84 = 7'h4e == _GEN_793 ? L0Memory_78 : _GEN_83; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_85 = 7'h4f == _GEN_793 ? L0Memory_79 : _GEN_84; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_86 = 7'h50 == _GEN_793 ? L0Memory_80 : _GEN_85; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_87 = 7'h51 == _GEN_793 ? L0Memory_81 : _GEN_86; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_88 = 7'h52 == _GEN_793 ? L0Memory_82 : _GEN_87; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_89 = 7'h53 == _GEN_793 ? L0Memory_83 : _GEN_88; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_90 = 7'h54 == _GEN_793 ? L0Memory_84 : _GEN_89; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_91 = 7'h55 == _GEN_793 ? L0Memory_85 : _GEN_90; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_92 = 7'h56 == _GEN_793 ? L0Memory_86 : _GEN_91; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_93 = 7'h57 == _GEN_793 ? L0Memory_87 : _GEN_92; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_94 = 7'h58 == _GEN_793 ? L0Memory_88 : _GEN_93; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_95 = 7'h59 == _GEN_793 ? L0Memory_89 : _GEN_94; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_96 = 7'h5a == _GEN_793 ? L0Memory_90 : _GEN_95; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_97 = 7'h5b == _GEN_793 ? L0Memory_91 : _GEN_96; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_98 = 7'h5c == _GEN_793 ? L0Memory_92 : _GEN_97; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_99 = 7'h5d == _GEN_793 ? L0Memory_93 : _GEN_98; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_100 = 7'h5e == _GEN_793 ? L0Memory_94 : _GEN_99; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_101 = 7'h5f == _GEN_793 ? L0Memory_95 : _GEN_100; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_102 = 7'h60 == _GEN_793 ? L0Memory_96 : _GEN_101; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_103 = 7'h61 == _GEN_793 ? L0Memory_97 : _GEN_102; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_104 = 7'h62 == _GEN_793 ? L0Memory_98 : _GEN_103; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_105 = 7'h63 == _GEN_793 ? L0Memory_99 : _GEN_104; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire  _GEN_575 = _T_12 ? 1'h0 : _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 157:12]
  wire  sel5 = _T_3 ? 1'h0 : _GEN_575; // @[Conditional.scala 40:58 PEArray.scala 112:12]
  reg [15:0] mux2out_reg; // @[PEArray.scala 90:28]
  reg [15:0] mux3out_reg; // @[PEArray.scala 91:28]
  reg [9:0] count; // @[PEArray.scala 101:22]
  reg [5:0] GRU_out_width; // @[PEArray.scala 104:26]
  wire [7:0] _GEN_118 = io_control_signal_mask[1] ? 8'h0 : {{2'd0}, GRU_out_width}; // @[PEArray.scala 116:57 PEArray.scala 145:23 PEArray.scala 104:26]
  wire [9:0] _count_T_1 = count + 10'h1; // @[PEArray.scala 162:24]
  wire [9:0] _GEN_120 = count != 10'h33 ? _count_T_1 : count; // @[PEArray.scala 161:27 PEArray.scala 162:15 PEArray.scala 101:22]
  wire [9:0] _GEN_124 = count != 10'h188 ? _count_T_1 : count; // @[PEArray.scala 183:28 PEArray.scala 184:15 PEArray.scala 101:22]
  wire [9:0] _GEN_125 = count == 10'h188 ? 10'h0 : _GEN_124; // @[PEArray.scala 186:28 PEArray.scala 187:15]
  wire [2:0] _GEN_126 = count == 10'h188 ? 3'h0 : state; // @[PEArray.scala 186:28 PEArray.scala 188:15 PEArray.scala 100:22]
  wire [9:0] _GEN_127 = count != 10'h0 ? _count_T_1 : count; // @[PEArray.scala 192:32 PEArray.scala 193:15 PEArray.scala 101:22]
  wire  _T_24 = count == 10'h0; // @[PEArray.scala 195:18]
  wire [5:0] _GEN_128 = count == 10'h0 ? 6'h0 : L0Index; // @[PEArray.scala 195:26 PEArray.scala 196:17 PEArray.scala 39:24]
  wire [9:0] _T_27 = 10'h0 - 10'h1; // @[PEArray.scala 198:51]
  wire [15:0] _GEN_129 = 6'h0 == L0Index ? io_FromL1 : L0Memory_0; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_130 = 6'h1 == L0Index ? io_FromL1 : L0Memory_1; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_131 = 6'h2 == L0Index ? io_FromL1 : L0Memory_2; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_132 = 6'h3 == L0Index ? io_FromL1 : L0Memory_3; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_133 = 6'h4 == L0Index ? io_FromL1 : L0Memory_4; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_134 = 6'h5 == L0Index ? io_FromL1 : L0Memory_5; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_135 = 6'h6 == L0Index ? io_FromL1 : L0Memory_6; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_136 = 6'h7 == L0Index ? io_FromL1 : L0Memory_7; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_137 = 6'h8 == L0Index ? io_FromL1 : L0Memory_8; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_138 = 6'h9 == L0Index ? io_FromL1 : L0Memory_9; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_139 = 6'ha == L0Index ? io_FromL1 : L0Memory_10; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_140 = 6'hb == L0Index ? io_FromL1 : L0Memory_11; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_141 = 6'hc == L0Index ? io_FromL1 : L0Memory_12; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_142 = 6'hd == L0Index ? io_FromL1 : L0Memory_13; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_143 = 6'he == L0Index ? io_FromL1 : L0Memory_14; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_144 = 6'hf == L0Index ? io_FromL1 : L0Memory_15; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_145 = 6'h10 == L0Index ? io_FromL1 : L0Memory_16; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_146 = 6'h11 == L0Index ? io_FromL1 : L0Memory_17; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_147 = 6'h12 == L0Index ? io_FromL1 : L0Memory_18; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_148 = 6'h13 == L0Index ? io_FromL1 : L0Memory_19; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_149 = 6'h14 == L0Index ? io_FromL1 : L0Memory_20; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_150 = 6'h15 == L0Index ? io_FromL1 : L0Memory_21; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_151 = 6'h16 == L0Index ? io_FromL1 : L0Memory_22; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_152 = 6'h17 == L0Index ? io_FromL1 : L0Memory_23; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_153 = 6'h18 == L0Index ? io_FromL1 : L0Memory_24; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_154 = 6'h19 == L0Index ? io_FromL1 : L0Memory_25; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_155 = 6'h1a == L0Index ? io_FromL1 : L0Memory_26; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_156 = 6'h1b == L0Index ? io_FromL1 : L0Memory_27; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_157 = 6'h1c == L0Index ? io_FromL1 : L0Memory_28; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_158 = 6'h1d == L0Index ? io_FromL1 : L0Memory_29; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_159 = 6'h1e == L0Index ? io_FromL1 : L0Memory_30; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_160 = 6'h1f == L0Index ? io_FromL1 : L0Memory_31; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_161 = 6'h20 == L0Index ? io_FromL1 : L0Memory_32; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_162 = 6'h21 == L0Index ? io_FromL1 : L0Memory_33; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_163 = 6'h22 == L0Index ? io_FromL1 : L0Memory_34; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_164 = 6'h23 == L0Index ? io_FromL1 : L0Memory_35; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_165 = 6'h24 == L0Index ? io_FromL1 : L0Memory_36; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_166 = 6'h25 == L0Index ? io_FromL1 : L0Memory_37; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_167 = 6'h26 == L0Index ? io_FromL1 : L0Memory_38; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_168 = 6'h27 == L0Index ? io_FromL1 : L0Memory_39; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_169 = 6'h28 == L0Index ? io_FromL1 : L0Memory_40; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_170 = 6'h29 == L0Index ? io_FromL1 : L0Memory_41; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_171 = 6'h2a == L0Index ? io_FromL1 : L0Memory_42; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_172 = 6'h2b == L0Index ? io_FromL1 : L0Memory_43; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_173 = 6'h2c == L0Index ? io_FromL1 : L0Memory_44; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_174 = 6'h2d == L0Index ? io_FromL1 : L0Memory_45; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_175 = 6'h2e == L0Index ? io_FromL1 : L0Memory_46; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_176 = 6'h2f == L0Index ? io_FromL1 : L0Memory_47; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_177 = 6'h30 == L0Index ? io_FromL1 : L0Memory_48; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_178 = 6'h31 == L0Index ? io_FromL1 : L0Memory_49; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_179 = 6'h32 == L0Index ? io_FromL1 : L0Memory_50; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_180 = 6'h33 == L0Index ? io_FromL1 : L0Memory_51; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_181 = 6'h34 == L0Index ? io_FromL1 : L0Memory_52; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_182 = 6'h35 == L0Index ? io_FromL1 : L0Memory_53; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_183 = 6'h36 == L0Index ? io_FromL1 : L0Memory_54; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_184 = 6'h37 == L0Index ? io_FromL1 : L0Memory_55; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_185 = 6'h38 == L0Index ? io_FromL1 : L0Memory_56; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_186 = 6'h39 == L0Index ? io_FromL1 : L0Memory_57; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_187 = 6'h3a == L0Index ? io_FromL1 : L0Memory_58; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_188 = 6'h3b == L0Index ? io_FromL1 : L0Memory_59; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_189 = 6'h3c == L0Index ? io_FromL1 : L0Memory_60; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_190 = 6'h3d == L0Index ? io_FromL1 : L0Memory_61; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_191 = 6'h3e == L0Index ? io_FromL1 : L0Memory_62; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_192 = 6'h3f == L0Index ? io_FromL1 : L0Memory_63; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_193 = 7'h40 == _GEN_793 ? io_FromL1 : L0Memory_64; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_194 = 7'h41 == _GEN_793 ? io_FromL1 : L0Memory_65; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_195 = 7'h42 == _GEN_793 ? io_FromL1 : L0Memory_66; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_196 = 7'h43 == _GEN_793 ? io_FromL1 : L0Memory_67; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_197 = 7'h44 == _GEN_793 ? io_FromL1 : L0Memory_68; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_198 = 7'h45 == _GEN_793 ? io_FromL1 : L0Memory_69; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_199 = 7'h46 == _GEN_793 ? io_FromL1 : L0Memory_70; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_200 = 7'h47 == _GEN_793 ? io_FromL1 : L0Memory_71; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_201 = 7'h48 == _GEN_793 ? io_FromL1 : L0Memory_72; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_202 = 7'h49 == _GEN_793 ? io_FromL1 : L0Memory_73; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_203 = 7'h4a == _GEN_793 ? io_FromL1 : L0Memory_74; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_204 = 7'h4b == _GEN_793 ? io_FromL1 : L0Memory_75; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_205 = 7'h4c == _GEN_793 ? io_FromL1 : L0Memory_76; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_206 = 7'h4d == _GEN_793 ? io_FromL1 : L0Memory_77; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_207 = 7'h4e == _GEN_793 ? io_FromL1 : L0Memory_78; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_208 = 7'h4f == _GEN_793 ? io_FromL1 : L0Memory_79; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_209 = 7'h50 == _GEN_793 ? io_FromL1 : L0Memory_80; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_210 = 7'h51 == _GEN_793 ? io_FromL1 : L0Memory_81; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_211 = 7'h52 == _GEN_793 ? io_FromL1 : L0Memory_82; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_212 = 7'h53 == _GEN_793 ? io_FromL1 : L0Memory_83; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_213 = 7'h54 == _GEN_793 ? io_FromL1 : L0Memory_84; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_214 = 7'h55 == _GEN_793 ? io_FromL1 : L0Memory_85; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_215 = 7'h56 == _GEN_793 ? io_FromL1 : L0Memory_86; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_216 = 7'h57 == _GEN_793 ? io_FromL1 : L0Memory_87; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_217 = 7'h58 == _GEN_793 ? io_FromL1 : L0Memory_88; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_218 = 7'h59 == _GEN_793 ? io_FromL1 : L0Memory_89; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_219 = 7'h5a == _GEN_793 ? io_FromL1 : L0Memory_90; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_220 = 7'h5b == _GEN_793 ? io_FromL1 : L0Memory_91; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_221 = 7'h5c == _GEN_793 ? io_FromL1 : L0Memory_92; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_222 = 7'h5d == _GEN_793 ? io_FromL1 : L0Memory_93; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_223 = 7'h5e == _GEN_793 ? io_FromL1 : L0Memory_94; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_224 = 7'h5f == _GEN_793 ? io_FromL1 : L0Memory_95; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_225 = 7'h60 == _GEN_793 ? io_FromL1 : L0Memory_96; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_226 = 7'h61 == _GEN_793 ? io_FromL1 : L0Memory_97; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_227 = 7'h62 == _GEN_793 ? io_FromL1 : L0Memory_98; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_228 = 7'h63 == _GEN_793 ? io_FromL1 : L0Memory_99; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [5:0] _L0Index_T_2 = L0Index + 6'h1; // @[PEArray.scala 200:28]
  wire [15:0] _GEN_229 = count >= 10'h1 & count <= _T_27 ? _GEN_129 : L0Memory_0; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_230 = count >= 10'h1 & count <= _T_27 ? _GEN_130 : L0Memory_1; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_231 = count >= 10'h1 & count <= _T_27 ? _GEN_131 : L0Memory_2; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_232 = count >= 10'h1 & count <= _T_27 ? _GEN_132 : L0Memory_3; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_233 = count >= 10'h1 & count <= _T_27 ? _GEN_133 : L0Memory_4; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_234 = count >= 10'h1 & count <= _T_27 ? _GEN_134 : L0Memory_5; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_235 = count >= 10'h1 & count <= _T_27 ? _GEN_135 : L0Memory_6; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_236 = count >= 10'h1 & count <= _T_27 ? _GEN_136 : L0Memory_7; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_237 = count >= 10'h1 & count <= _T_27 ? _GEN_137 : L0Memory_8; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_238 = count >= 10'h1 & count <= _T_27 ? _GEN_138 : L0Memory_9; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_239 = count >= 10'h1 & count <= _T_27 ? _GEN_139 : L0Memory_10; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_240 = count >= 10'h1 & count <= _T_27 ? _GEN_140 : L0Memory_11; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_241 = count >= 10'h1 & count <= _T_27 ? _GEN_141 : L0Memory_12; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_242 = count >= 10'h1 & count <= _T_27 ? _GEN_142 : L0Memory_13; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_243 = count >= 10'h1 & count <= _T_27 ? _GEN_143 : L0Memory_14; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_244 = count >= 10'h1 & count <= _T_27 ? _GEN_144 : L0Memory_15; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_245 = count >= 10'h1 & count <= _T_27 ? _GEN_145 : L0Memory_16; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_246 = count >= 10'h1 & count <= _T_27 ? _GEN_146 : L0Memory_17; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_247 = count >= 10'h1 & count <= _T_27 ? _GEN_147 : L0Memory_18; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_248 = count >= 10'h1 & count <= _T_27 ? _GEN_148 : L0Memory_19; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_249 = count >= 10'h1 & count <= _T_27 ? _GEN_149 : L0Memory_20; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_250 = count >= 10'h1 & count <= _T_27 ? _GEN_150 : L0Memory_21; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_251 = count >= 10'h1 & count <= _T_27 ? _GEN_151 : L0Memory_22; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_252 = count >= 10'h1 & count <= _T_27 ? _GEN_152 : L0Memory_23; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_253 = count >= 10'h1 & count <= _T_27 ? _GEN_153 : L0Memory_24; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_254 = count >= 10'h1 & count <= _T_27 ? _GEN_154 : L0Memory_25; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_255 = count >= 10'h1 & count <= _T_27 ? _GEN_155 : L0Memory_26; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_256 = count >= 10'h1 & count <= _T_27 ? _GEN_156 : L0Memory_27; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_257 = count >= 10'h1 & count <= _T_27 ? _GEN_157 : L0Memory_28; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_258 = count >= 10'h1 & count <= _T_27 ? _GEN_158 : L0Memory_29; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_259 = count >= 10'h1 & count <= _T_27 ? _GEN_159 : L0Memory_30; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_260 = count >= 10'h1 & count <= _T_27 ? _GEN_160 : L0Memory_31; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_261 = count >= 10'h1 & count <= _T_27 ? _GEN_161 : L0Memory_32; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_262 = count >= 10'h1 & count <= _T_27 ? _GEN_162 : L0Memory_33; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_263 = count >= 10'h1 & count <= _T_27 ? _GEN_163 : L0Memory_34; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_264 = count >= 10'h1 & count <= _T_27 ? _GEN_164 : L0Memory_35; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_265 = count >= 10'h1 & count <= _T_27 ? _GEN_165 : L0Memory_36; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_266 = count >= 10'h1 & count <= _T_27 ? _GEN_166 : L0Memory_37; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_267 = count >= 10'h1 & count <= _T_27 ? _GEN_167 : L0Memory_38; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_268 = count >= 10'h1 & count <= _T_27 ? _GEN_168 : L0Memory_39; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_269 = count >= 10'h1 & count <= _T_27 ? _GEN_169 : L0Memory_40; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_270 = count >= 10'h1 & count <= _T_27 ? _GEN_170 : L0Memory_41; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_271 = count >= 10'h1 & count <= _T_27 ? _GEN_171 : L0Memory_42; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_272 = count >= 10'h1 & count <= _T_27 ? _GEN_172 : L0Memory_43; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_273 = count >= 10'h1 & count <= _T_27 ? _GEN_173 : L0Memory_44; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_274 = count >= 10'h1 & count <= _T_27 ? _GEN_174 : L0Memory_45; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_275 = count >= 10'h1 & count <= _T_27 ? _GEN_175 : L0Memory_46; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_276 = count >= 10'h1 & count <= _T_27 ? _GEN_176 : L0Memory_47; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_277 = count >= 10'h1 & count <= _T_27 ? _GEN_177 : L0Memory_48; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_278 = count >= 10'h1 & count <= _T_27 ? _GEN_178 : L0Memory_49; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_279 = count >= 10'h1 & count <= _T_27 ? _GEN_179 : L0Memory_50; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_280 = count >= 10'h1 & count <= _T_27 ? _GEN_180 : L0Memory_51; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_281 = count >= 10'h1 & count <= _T_27 ? _GEN_181 : L0Memory_52; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_282 = count >= 10'h1 & count <= _T_27 ? _GEN_182 : L0Memory_53; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_283 = count >= 10'h1 & count <= _T_27 ? _GEN_183 : L0Memory_54; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_284 = count >= 10'h1 & count <= _T_27 ? _GEN_184 : L0Memory_55; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_285 = count >= 10'h1 & count <= _T_27 ? _GEN_185 : L0Memory_56; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_286 = count >= 10'h1 & count <= _T_27 ? _GEN_186 : L0Memory_57; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_287 = count >= 10'h1 & count <= _T_27 ? _GEN_187 : L0Memory_58; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_288 = count >= 10'h1 & count <= _T_27 ? _GEN_188 : L0Memory_59; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_289 = count >= 10'h1 & count <= _T_27 ? _GEN_189 : L0Memory_60; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_290 = count >= 10'h1 & count <= _T_27 ? _GEN_190 : L0Memory_61; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_291 = count >= 10'h1 & count <= _T_27 ? _GEN_191 : L0Memory_62; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_292 = count >= 10'h1 & count <= _T_27 ? _GEN_192 : L0Memory_63; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_293 = count >= 10'h1 & count <= _T_27 ? _GEN_193 : L0Memory_64; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_294 = count >= 10'h1 & count <= _T_27 ? _GEN_194 : L0Memory_65; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_295 = count >= 10'h1 & count <= _T_27 ? _GEN_195 : L0Memory_66; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_296 = count >= 10'h1 & count <= _T_27 ? _GEN_196 : L0Memory_67; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_297 = count >= 10'h1 & count <= _T_27 ? _GEN_197 : L0Memory_68; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_298 = count >= 10'h1 & count <= _T_27 ? _GEN_198 : L0Memory_69; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_299 = count >= 10'h1 & count <= _T_27 ? _GEN_199 : L0Memory_70; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_300 = count >= 10'h1 & count <= _T_27 ? _GEN_200 : L0Memory_71; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_301 = count >= 10'h1 & count <= _T_27 ? _GEN_201 : L0Memory_72; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_302 = count >= 10'h1 & count <= _T_27 ? _GEN_202 : L0Memory_73; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_303 = count >= 10'h1 & count <= _T_27 ? _GEN_203 : L0Memory_74; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_304 = count >= 10'h1 & count <= _T_27 ? _GEN_204 : L0Memory_75; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_305 = count >= 10'h1 & count <= _T_27 ? _GEN_205 : L0Memory_76; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_306 = count >= 10'h1 & count <= _T_27 ? _GEN_206 : L0Memory_77; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_307 = count >= 10'h1 & count <= _T_27 ? _GEN_207 : L0Memory_78; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_308 = count >= 10'h1 & count <= _T_27 ? _GEN_208 : L0Memory_79; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_309 = count >= 10'h1 & count <= _T_27 ? _GEN_209 : L0Memory_80; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_310 = count >= 10'h1 & count <= _T_27 ? _GEN_210 : L0Memory_81; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_311 = count >= 10'h1 & count <= _T_27 ? _GEN_211 : L0Memory_82; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_312 = count >= 10'h1 & count <= _T_27 ? _GEN_212 : L0Memory_83; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_313 = count >= 10'h1 & count <= _T_27 ? _GEN_213 : L0Memory_84; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_314 = count >= 10'h1 & count <= _T_27 ? _GEN_214 : L0Memory_85; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_315 = count >= 10'h1 & count <= _T_27 ? _GEN_215 : L0Memory_86; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_316 = count >= 10'h1 & count <= _T_27 ? _GEN_216 : L0Memory_87; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_317 = count >= 10'h1 & count <= _T_27 ? _GEN_217 : L0Memory_88; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_318 = count >= 10'h1 & count <= _T_27 ? _GEN_218 : L0Memory_89; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_319 = count >= 10'h1 & count <= _T_27 ? _GEN_219 : L0Memory_90; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_320 = count >= 10'h1 & count <= _T_27 ? _GEN_220 : L0Memory_91; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_321 = count >= 10'h1 & count <= _T_27 ? _GEN_221 : L0Memory_92; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_322 = count >= 10'h1 & count <= _T_27 ? _GEN_222 : L0Memory_93; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_323 = count >= 10'h1 & count <= _T_27 ? _GEN_223 : L0Memory_94; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_324 = count >= 10'h1 & count <= _T_27 ? _GEN_224 : L0Memory_95; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_325 = count >= 10'h1 & count <= _T_27 ? _GEN_225 : L0Memory_96; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_326 = count >= 10'h1 & count <= _T_27 ? _GEN_226 : L0Memory_97; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_327 = count >= 10'h1 & count <= _T_27 ? _GEN_227 : L0Memory_98; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_328 = count >= 10'h1 & count <= _T_27 ? _GEN_228 : L0Memory_99; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [5:0] _GEN_329 = count >= 10'h1 & count <= _T_27 ? _L0Index_T_2 : _GEN_128; // @[PEArray.scala 198:59 PEArray.scala 200:17]
  wire [9:0] _GEN_330 = _T_24 ? 10'h0 : _GEN_127; // @[PEArray.scala 202:32 PEArray.scala 203:15]
  wire [2:0] _GEN_331 = _T_24 ? 3'h0 : state; // @[PEArray.scala 202:32 PEArray.scala 204:15 PEArray.scala 100:22]
  wire [9:0] _GEN_865 = {{4'd0}, GRU_out_width}; // @[PEArray.scala 220:19]
  wire [9:0] _GEN_0 = count % _GEN_865; // @[PEArray.scala 220:19]
  wire [5:0] _T_36 = _GEN_0[5:0]; // @[PEArray.scala 220:19]
  wire [5:0] _T_38 = GRU_out_width - 6'h1; // @[PEArray.scala 220:55]
  wire [5:0] _GEN_334 = _T_36 == _T_38 ? _L0Index_T_2 : 6'h0; // @[PEArray.scala 220:62 PEArray.scala 221:17 PEArray.scala 214:15]
  wire [5:0] _GEN_346 = _T_41 ? _GEN_334 : L0Index; // @[Conditional.scala 39:67 PEArray.scala 39:24]
  wire [9:0] _GEN_347 = _T_41 ? _GEN_330 : count; // @[Conditional.scala 39:67 PEArray.scala 101:22]
  wire [2:0] _GEN_348 = _T_41 ? _GEN_331 : state; // @[Conditional.scala 39:67 PEArray.scala 100:22]
  wire [5:0] _GEN_353 = _T_31 ? _GEN_334 : _GEN_346; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_354 = _T_31 ? _GEN_330 : _GEN_347; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_355 = _T_31 ? _GEN_331 : _GEN_348; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_356 = _T_22 ? _GEN_330 : _GEN_354; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_357 = _T_22 ? _GEN_329 : _GEN_353; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_458 = _T_22 ? _GEN_331 : _GEN_355; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_690 = _T_3 ? _GEN_118 : {{2'd0}, GRU_out_width}; // @[Conditional.scala 40:58 PEArray.scala 104:26]
  FP16MulAdder FP16MAC ( // @[PEArray.scala 72:23]
    .io_a(FP16MAC_io_a),
    .io_b(FP16MAC_io_b),
    .io_c(FP16MAC_io_c),
    .io_out(FP16MAC_io_out)
  );
  assign io_ToRightPE = mux3out_reg; // @[PEArray.scala 95:16]
  assign io_ToBelowPE = mux2out_reg; // @[PEArray.scala 94:16]
  assign FP16MAC_io_a = sel1 ? io_FromL1 : io_FromLeftPE; // @[PEArray.scala 50:14 PEArray.scala 50:23 PEArray.scala 51:24]
  assign FP16MAC_io_b = sel5 ? mux4out : _GEN_105; // @[PEArray.scala 77:13 PEArray.scala 78:18 PEArray.scala 81:18]
  assign FP16MAC_io_c = sel5 ? _GEN_105 : mux4out; // @[PEArray.scala 77:13 PEArray.scala 79:18 PEArray.scala 82:18]
  always @(posedge clock) begin
    if (reset) begin // @[PEArray.scala 39:24]
      L0Index <= 6'h0; // @[PEArray.scala 39:24]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h1; // @[PEArray.scala 159:15]
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        L0Index <= 6'hd; // @[PEArray.scala 181:15]
      end else begin
        L0Index <= _GEN_357;
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_0 <= _GEN_229;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_1 <= _GEN_230;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_2 <= _GEN_231;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_3 <= _GEN_232;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_4 <= _GEN_233;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_5 <= _GEN_234;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_6 <= _GEN_235;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_7 <= _GEN_236;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_8 <= _GEN_237;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_9 <= _GEN_238;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_10 <= _GEN_239;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_11 <= _GEN_240;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_12 <= _GEN_241;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_13 <= _GEN_242;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_14 <= _GEN_243;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_15 <= _GEN_244;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_16 <= _GEN_245;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_17 <= _GEN_246;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_18 <= _GEN_247;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_19 <= _GEN_248;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_20 <= _GEN_249;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_21 <= _GEN_250;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_22 <= _GEN_251;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_23 <= _GEN_252;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_24 <= _GEN_253;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_25 <= _GEN_254;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_26 <= _GEN_255;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_27 <= _GEN_256;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_28 <= _GEN_257;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_29 <= _GEN_258;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_30 <= _GEN_259;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_31 <= _GEN_260;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_32 <= _GEN_261;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_33 <= _GEN_262;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_34 <= _GEN_263;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_35 <= _GEN_264;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_36 <= _GEN_265;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_37 <= _GEN_266;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_38 <= _GEN_267;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_39 <= _GEN_268;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_40 <= _GEN_269;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_41 <= _GEN_270;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_42 <= _GEN_271;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_43 <= _GEN_272;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_44 <= _GEN_273;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_45 <= _GEN_274;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_46 <= _GEN_275;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_47 <= _GEN_276;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_48 <= _GEN_277;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_49 <= _GEN_278;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_50 <= _GEN_279;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_51 <= _GEN_280;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_52 <= _GEN_281;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_53 <= _GEN_282;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_54 <= _GEN_283;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_55 <= _GEN_284;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_56 <= _GEN_285;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_57 <= _GEN_286;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_58 <= _GEN_287;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_59 <= _GEN_288;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_60 <= _GEN_289;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_61 <= _GEN_290;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_62 <= _GEN_291;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_63 <= _GEN_292;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_64 <= _GEN_293;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_65 <= _GEN_294;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_66 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_67 <= _GEN_296;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_68 <= _GEN_297;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_69 <= _GEN_298;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_70 <= _GEN_299;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_71 <= _GEN_300;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_72 <= _GEN_301;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_73 <= _GEN_302;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_74 <= _GEN_303;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_75 <= _GEN_304;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_76 <= _GEN_305;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_77 <= _GEN_306;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_78 <= _GEN_307;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_79 <= _GEN_308;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_80 <= _GEN_309;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_81 <= _GEN_310;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_82 <= _GEN_311;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_83 <= _GEN_312;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_84 <= _GEN_313;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_85 <= _GEN_314;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_86 <= _GEN_315;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_87 <= _GEN_316;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_88 <= _GEN_317;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_89 <= _GEN_318;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_90 <= _GEN_319;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_91 <= _GEN_320;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_92 <= _GEN_321;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_93 <= _GEN_322;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_94 <= _GEN_323;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_95 <= _GEN_324;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_96 <= _GEN_325;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_97 <= _GEN_326;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_98 <= _GEN_327;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_99 <= _GEN_328;
          end
        end
      end
    end
    if (reset) begin // @[PEArray.scala 100:22]
      state <= 3'h0; // @[PEArray.scala 100:22]
    end else if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[1]) begin // @[PEArray.scala 116:57]
        state <= 3'h1;
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      if (count == 10'h33) begin // @[PEArray.scala 164:27]
        state <= 3'h0; // @[PEArray.scala 166:15]
      end
    end else if (_T_16) begin // @[Conditional.scala 39:67]
      state <= _GEN_126;
    end else begin
      state <= _GEN_458;
    end
    if (reset) begin // @[PEArray.scala 90:28]
      mux2out_reg <= 16'h0; // @[PEArray.scala 90:28]
    end else begin
      mux2out_reg <= MAC_out; // @[PEArray.scala 90:28]
    end
    if (reset) begin // @[PEArray.scala 91:28]
      mux3out_reg <= 16'h0; // @[PEArray.scala 91:28]
    end else if (sel3) begin // @[PEArray.scala 56:14]
      mux3out_reg <= MAC_out; // @[PEArray.scala 56:23]
    end else if (sel1) begin // @[PEArray.scala 50:14]
      mux3out_reg <= io_FromL1; // @[PEArray.scala 50:23]
    end else begin
      mux3out_reg <= io_FromLeftPE; // @[PEArray.scala 51:24]
    end
    if (reset) begin // @[PEArray.scala 101:22]
      count <= 10'h0; // @[PEArray.scala 101:22]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        if (count == 10'h33) begin // @[PEArray.scala 164:27]
          count <= 10'h0; // @[PEArray.scala 165:15]
        end else begin
          count <= _GEN_120;
        end
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        count <= _GEN_125;
      end else begin
        count <= _GEN_356;
      end
    end
    GRU_out_width <= _GEN_690[5:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  L0Index = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  L0Memory_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  L0Memory_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  L0Memory_2 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  L0Memory_3 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  L0Memory_4 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  L0Memory_5 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  L0Memory_6 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  L0Memory_7 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  L0Memory_8 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  L0Memory_9 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  L0Memory_10 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  L0Memory_11 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  L0Memory_12 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  L0Memory_13 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  L0Memory_14 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  L0Memory_15 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  L0Memory_16 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  L0Memory_17 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  L0Memory_18 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  L0Memory_19 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  L0Memory_20 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  L0Memory_21 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  L0Memory_22 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  L0Memory_23 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  L0Memory_24 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  L0Memory_25 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  L0Memory_26 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  L0Memory_27 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  L0Memory_28 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  L0Memory_29 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  L0Memory_30 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  L0Memory_31 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  L0Memory_32 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  L0Memory_33 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  L0Memory_34 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  L0Memory_35 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  L0Memory_36 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  L0Memory_37 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  L0Memory_38 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  L0Memory_39 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  L0Memory_40 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  L0Memory_41 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  L0Memory_42 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  L0Memory_43 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  L0Memory_44 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  L0Memory_45 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  L0Memory_46 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  L0Memory_47 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  L0Memory_48 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  L0Memory_49 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  L0Memory_50 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  L0Memory_51 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  L0Memory_52 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  L0Memory_53 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  L0Memory_54 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  L0Memory_55 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  L0Memory_56 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  L0Memory_57 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  L0Memory_58 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  L0Memory_59 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  L0Memory_60 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  L0Memory_61 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  L0Memory_62 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  L0Memory_63 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  L0Memory_64 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  L0Memory_65 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  L0Memory_66 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  L0Memory_67 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  L0Memory_68 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  L0Memory_69 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  L0Memory_70 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  L0Memory_71 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  L0Memory_72 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  L0Memory_73 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  L0Memory_74 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  L0Memory_75 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  L0Memory_76 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  L0Memory_77 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  L0Memory_78 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  L0Memory_79 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  L0Memory_80 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  L0Memory_81 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  L0Memory_82 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  L0Memory_83 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  L0Memory_84 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  L0Memory_85 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  L0Memory_86 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  L0Memory_87 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  L0Memory_88 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  L0Memory_89 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  L0Memory_90 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  L0Memory_91 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  L0Memory_92 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  L0Memory_93 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  L0Memory_94 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  L0Memory_95 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  L0Memory_96 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  L0Memory_97 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  L0Memory_98 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  L0Memory_99 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  state = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  mux2out_reg = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  mux3out_reg = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  count = _RAND_104[9:0];
  _RAND_105 = {1{`RANDOM}};
  GRU_out_width = _RAND_105[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PE_32(
  input         clock,
  input         reset,
  input  [15:0] io_FromAbovePE,
  input  [15:0] io_FromLeftPE,
  input  [15:0] io_FromL1,
  input  [2:0]  io_control_signal_control,
  input  [9:0]  io_control_signal_count,
  input  [5:0]  io_control_signal_L0index,
  input  [11:0] io_control_signal_mask,
  input  [7:0]  io_control_signal_gru_out_width,
  output [15:0] io_ToRightPE,
  output [15:0] io_ToBelowPE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] FP16MAC_io_a; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_b; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_c; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_out; // @[PEArray.scala 72:23]
  reg [5:0] L0Index; // @[PEArray.scala 39:24]
  reg [15:0] L0Memory_0; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_1; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_2; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_3; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_4; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_5; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_6; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_7; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_8; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_9; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_10; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_11; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_12; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_13; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_14; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_15; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_16; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_17; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_18; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_19; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_20; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_21; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_22; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_23; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_24; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_25; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_26; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_27; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_28; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_29; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_30; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_31; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_32; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_33; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_34; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_35; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_36; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_37; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_38; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_39; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_40; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_41; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_42; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_43; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_44; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_45; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_46; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_47; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_48; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_49; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_50; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_51; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_52; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_53; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_54; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_55; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_56; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_57; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_58; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_59; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_60; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_61; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_62; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_63; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_64; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_65; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_66; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_67; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_68; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_69; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_70; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_71; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_72; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_73; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_74; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_75; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_76; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_77; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_78; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_79; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_80; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_81; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_82; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_83; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_84; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_85; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_86; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_87; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_88; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_89; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_90; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_91; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_92; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_93; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_94; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_95; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_96; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_97; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_98; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_99; // @[PEArray.scala 40:21]
  reg [2:0] state; // @[PEArray.scala 100:22]
  wire  _T_3 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_12 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_16 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_22 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_31 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_41 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_342 = _T_41 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 231:12 PEArray.scala 32:8]
  wire  _GEN_349 = _T_31 ? 1'h0 : _GEN_342; // @[Conditional.scala 39:67 PEArray.scala 208:12]
  wire  _GEN_459 = _T_22 | _GEN_349; // @[Conditional.scala 39:67 PEArray.scala 32:8]
  wire  _GEN_463 = _T_16 ? 1'h0 : _GEN_459; // @[Conditional.scala 39:67]
  wire  _GEN_572 = _T_12 | _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 149:12]
  wire  sel1 = _T_3 | _GEN_572; // @[Conditional.scala 40:58 PEArray.scala 108:12]
  wire [15:0] MAC_out = FP16MAC_io_out; // @[PEArray.scala 47:21 PEArray.scala 85:11]
  wire  _GEN_465 = _T_16 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 177:12]
  wire  _GEN_580 = _T_12 | _GEN_465; // @[Conditional.scala 39:67 PEArray.scala 34:8]
  wire  sel3 = _T_3 | _GEN_580; // @[Conditional.scala 40:58 PEArray.scala 110:12]
  wire [1:0] _GEN_344 = _T_41 ? 2'h2 : 2'h0; // @[Conditional.scala 39:67 PEArray.scala 233:12 PEArray.scala 35:8]
  wire [1:0] _GEN_351 = _T_31 ? 2'h2 : _GEN_344; // @[Conditional.scala 39:67 PEArray.scala 210:12]
  wire [1:0] _GEN_461 = _T_22 ? 2'h0 : _GEN_351; // @[Conditional.scala 39:67 PEArray.scala 35:8]
  wire [1:0] _GEN_466 = _T_16 ? 2'h0 : _GEN_461; // @[Conditional.scala 39:67 PEArray.scala 178:12]
  wire [1:0] _GEN_574 = _T_12 ? 2'h1 : _GEN_466; // @[Conditional.scala 39:67]
  wire [1:0] sel4 = _T_3 ? 2'h0 : _GEN_574; // @[Conditional.scala 40:58 PEArray.scala 111:12]
  wire [15:0] _GEN_3 = sel4 == 2'h2 ? io_FromL1 : 16'h0; // @[PEArray.scala 65:28 PEArray.scala 66:15 PEArray.scala 69:15]
  wire [15:0] _GEN_4 = sel4 == 2'h1 ? io_FromAbovePE : _GEN_3; // @[PEArray.scala 62:28 PEArray.scala 63:15]
  wire [15:0] mux4out = sel4 == 2'h0 ? 16'h0 : _GEN_4; // @[PEArray.scala 59:22 PEArray.scala 60:13]
  wire [15:0] _GEN_7 = 6'h1 == L0Index ? L0Memory_1 : L0Memory_0; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_8 = 6'h2 == L0Index ? L0Memory_2 : _GEN_7; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_9 = 6'h3 == L0Index ? L0Memory_3 : _GEN_8; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_10 = 6'h4 == L0Index ? L0Memory_4 : _GEN_9; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_11 = 6'h5 == L0Index ? L0Memory_5 : _GEN_10; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_12 = 6'h6 == L0Index ? L0Memory_6 : _GEN_11; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_13 = 6'h7 == L0Index ? L0Memory_7 : _GEN_12; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_14 = 6'h8 == L0Index ? L0Memory_8 : _GEN_13; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_15 = 6'h9 == L0Index ? L0Memory_9 : _GEN_14; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_16 = 6'ha == L0Index ? L0Memory_10 : _GEN_15; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_17 = 6'hb == L0Index ? L0Memory_11 : _GEN_16; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_18 = 6'hc == L0Index ? L0Memory_12 : _GEN_17; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_19 = 6'hd == L0Index ? L0Memory_13 : _GEN_18; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_20 = 6'he == L0Index ? L0Memory_14 : _GEN_19; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_21 = 6'hf == L0Index ? L0Memory_15 : _GEN_20; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_22 = 6'h10 == L0Index ? L0Memory_16 : _GEN_21; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_23 = 6'h11 == L0Index ? L0Memory_17 : _GEN_22; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_24 = 6'h12 == L0Index ? L0Memory_18 : _GEN_23; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_25 = 6'h13 == L0Index ? L0Memory_19 : _GEN_24; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_26 = 6'h14 == L0Index ? L0Memory_20 : _GEN_25; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_27 = 6'h15 == L0Index ? L0Memory_21 : _GEN_26; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_28 = 6'h16 == L0Index ? L0Memory_22 : _GEN_27; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_29 = 6'h17 == L0Index ? L0Memory_23 : _GEN_28; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_30 = 6'h18 == L0Index ? L0Memory_24 : _GEN_29; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_31 = 6'h19 == L0Index ? L0Memory_25 : _GEN_30; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_32 = 6'h1a == L0Index ? L0Memory_26 : _GEN_31; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_33 = 6'h1b == L0Index ? L0Memory_27 : _GEN_32; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_34 = 6'h1c == L0Index ? L0Memory_28 : _GEN_33; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_35 = 6'h1d == L0Index ? L0Memory_29 : _GEN_34; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_36 = 6'h1e == L0Index ? L0Memory_30 : _GEN_35; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_37 = 6'h1f == L0Index ? L0Memory_31 : _GEN_36; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_38 = 6'h20 == L0Index ? L0Memory_32 : _GEN_37; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_39 = 6'h21 == L0Index ? L0Memory_33 : _GEN_38; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_40 = 6'h22 == L0Index ? L0Memory_34 : _GEN_39; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_41 = 6'h23 == L0Index ? L0Memory_35 : _GEN_40; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_42 = 6'h24 == L0Index ? L0Memory_36 : _GEN_41; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_43 = 6'h25 == L0Index ? L0Memory_37 : _GEN_42; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_44 = 6'h26 == L0Index ? L0Memory_38 : _GEN_43; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_45 = 6'h27 == L0Index ? L0Memory_39 : _GEN_44; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_46 = 6'h28 == L0Index ? L0Memory_40 : _GEN_45; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_47 = 6'h29 == L0Index ? L0Memory_41 : _GEN_46; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_48 = 6'h2a == L0Index ? L0Memory_42 : _GEN_47; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_49 = 6'h2b == L0Index ? L0Memory_43 : _GEN_48; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_50 = 6'h2c == L0Index ? L0Memory_44 : _GEN_49; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_51 = 6'h2d == L0Index ? L0Memory_45 : _GEN_50; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_52 = 6'h2e == L0Index ? L0Memory_46 : _GEN_51; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_53 = 6'h2f == L0Index ? L0Memory_47 : _GEN_52; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_54 = 6'h30 == L0Index ? L0Memory_48 : _GEN_53; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_55 = 6'h31 == L0Index ? L0Memory_49 : _GEN_54; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_56 = 6'h32 == L0Index ? L0Memory_50 : _GEN_55; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_57 = 6'h33 == L0Index ? L0Memory_51 : _GEN_56; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_58 = 6'h34 == L0Index ? L0Memory_52 : _GEN_57; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_59 = 6'h35 == L0Index ? L0Memory_53 : _GEN_58; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_60 = 6'h36 == L0Index ? L0Memory_54 : _GEN_59; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_61 = 6'h37 == L0Index ? L0Memory_55 : _GEN_60; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_62 = 6'h38 == L0Index ? L0Memory_56 : _GEN_61; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_63 = 6'h39 == L0Index ? L0Memory_57 : _GEN_62; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_64 = 6'h3a == L0Index ? L0Memory_58 : _GEN_63; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_65 = 6'h3b == L0Index ? L0Memory_59 : _GEN_64; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_66 = 6'h3c == L0Index ? L0Memory_60 : _GEN_65; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_67 = 6'h3d == L0Index ? L0Memory_61 : _GEN_66; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_68 = 6'h3e == L0Index ? L0Memory_62 : _GEN_67; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_69 = 6'h3f == L0Index ? L0Memory_63 : _GEN_68; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [6:0] _GEN_793 = {{1'd0}, L0Index}; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_70 = 7'h40 == _GEN_793 ? L0Memory_64 : _GEN_69; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_71 = 7'h41 == _GEN_793 ? L0Memory_65 : _GEN_70; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_72 = 7'h42 == _GEN_793 ? L0Memory_66 : _GEN_71; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_73 = 7'h43 == _GEN_793 ? L0Memory_67 : _GEN_72; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_74 = 7'h44 == _GEN_793 ? L0Memory_68 : _GEN_73; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_75 = 7'h45 == _GEN_793 ? L0Memory_69 : _GEN_74; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_76 = 7'h46 == _GEN_793 ? L0Memory_70 : _GEN_75; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_77 = 7'h47 == _GEN_793 ? L0Memory_71 : _GEN_76; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_78 = 7'h48 == _GEN_793 ? L0Memory_72 : _GEN_77; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_79 = 7'h49 == _GEN_793 ? L0Memory_73 : _GEN_78; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_80 = 7'h4a == _GEN_793 ? L0Memory_74 : _GEN_79; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_81 = 7'h4b == _GEN_793 ? L0Memory_75 : _GEN_80; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_82 = 7'h4c == _GEN_793 ? L0Memory_76 : _GEN_81; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_83 = 7'h4d == _GEN_793 ? L0Memory_77 : _GEN_82; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_84 = 7'h4e == _GEN_793 ? L0Memory_78 : _GEN_83; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_85 = 7'h4f == _GEN_793 ? L0Memory_79 : _GEN_84; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_86 = 7'h50 == _GEN_793 ? L0Memory_80 : _GEN_85; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_87 = 7'h51 == _GEN_793 ? L0Memory_81 : _GEN_86; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_88 = 7'h52 == _GEN_793 ? L0Memory_82 : _GEN_87; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_89 = 7'h53 == _GEN_793 ? L0Memory_83 : _GEN_88; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_90 = 7'h54 == _GEN_793 ? L0Memory_84 : _GEN_89; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_91 = 7'h55 == _GEN_793 ? L0Memory_85 : _GEN_90; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_92 = 7'h56 == _GEN_793 ? L0Memory_86 : _GEN_91; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_93 = 7'h57 == _GEN_793 ? L0Memory_87 : _GEN_92; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_94 = 7'h58 == _GEN_793 ? L0Memory_88 : _GEN_93; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_95 = 7'h59 == _GEN_793 ? L0Memory_89 : _GEN_94; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_96 = 7'h5a == _GEN_793 ? L0Memory_90 : _GEN_95; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_97 = 7'h5b == _GEN_793 ? L0Memory_91 : _GEN_96; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_98 = 7'h5c == _GEN_793 ? L0Memory_92 : _GEN_97; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_99 = 7'h5d == _GEN_793 ? L0Memory_93 : _GEN_98; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_100 = 7'h5e == _GEN_793 ? L0Memory_94 : _GEN_99; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_101 = 7'h5f == _GEN_793 ? L0Memory_95 : _GEN_100; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_102 = 7'h60 == _GEN_793 ? L0Memory_96 : _GEN_101; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_103 = 7'h61 == _GEN_793 ? L0Memory_97 : _GEN_102; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_104 = 7'h62 == _GEN_793 ? L0Memory_98 : _GEN_103; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_105 = 7'h63 == _GEN_793 ? L0Memory_99 : _GEN_104; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire  _GEN_575 = _T_12 ? 1'h0 : _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 157:12]
  wire  sel5 = _T_3 ? 1'h0 : _GEN_575; // @[Conditional.scala 40:58 PEArray.scala 112:12]
  reg [15:0] mux2out_reg; // @[PEArray.scala 90:28]
  reg [15:0] mux3out_reg; // @[PEArray.scala 91:28]
  reg [9:0] count; // @[PEArray.scala 101:22]
  reg [9:0] count_max; // @[PEArray.scala 102:22]
  reg [5:0] L0index_begin; // @[PEArray.scala 103:26]
  reg [5:0] GRU_out_width; // @[PEArray.scala 104:26]
  wire  _T_6 = 3'h0 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_7 = 3'h1 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_8 = 3'h2 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_9 = 3'h3 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_10 = 3'h4 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_11 = 3'h5 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_109 = _T_11 ? 3'h5 : state; // @[Conditional.scala 39:67 PEArray.scala 140:19 PEArray.scala 100:22]
  wire [2:0] _GEN_110 = _T_10 ? 3'h4 : _GEN_109; // @[Conditional.scala 39:67 PEArray.scala 136:19]
  wire [2:0] _GEN_111 = _T_9 ? 3'h3 : _GEN_110; // @[Conditional.scala 39:67 PEArray.scala 132:19]
  wire [2:0] _GEN_112 = _T_8 ? 3'h2 : _GEN_111; // @[Conditional.scala 39:67 PEArray.scala 128:19]
  wire [2:0] _GEN_113 = _T_7 ? 3'h1 : _GEN_112; // @[Conditional.scala 39:67 PEArray.scala 124:19]
  wire [7:0] _GEN_118 = io_control_signal_mask[1] ? io_control_signal_gru_out_width : {{2'd0}, GRU_out_width}; // @[PEArray.scala 116:57 PEArray.scala 145:23 PEArray.scala 104:26]
  wire [9:0] _count_T_1 = count + 10'h1; // @[PEArray.scala 162:24]
  wire [9:0] _GEN_120 = count != 10'h33 ? _count_T_1 : count; // @[PEArray.scala 161:27 PEArray.scala 162:15 PEArray.scala 101:22]
  wire [9:0] _GEN_124 = count != 10'h188 ? _count_T_1 : count; // @[PEArray.scala 183:28 PEArray.scala 184:15 PEArray.scala 101:22]
  wire [9:0] _GEN_125 = count == 10'h188 ? 10'h0 : _GEN_124; // @[PEArray.scala 186:28 PEArray.scala 187:15]
  wire [2:0] _GEN_126 = count == 10'h188 ? 3'h0 : state; // @[PEArray.scala 186:28 PEArray.scala 188:15 PEArray.scala 100:22]
  wire [9:0] _GEN_127 = count != count_max ? _count_T_1 : count; // @[PEArray.scala 192:32 PEArray.scala 193:15 PEArray.scala 101:22]
  wire [5:0] _GEN_128 = count == 10'h0 ? L0index_begin : L0Index; // @[PEArray.scala 195:26 PEArray.scala 196:17 PEArray.scala 39:24]
  wire [9:0] _T_27 = count_max - 10'h1; // @[PEArray.scala 198:51]
  wire [15:0] _GEN_129 = 6'h0 == L0Index ? io_FromL1 : L0Memory_0; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_130 = 6'h1 == L0Index ? io_FromL1 : L0Memory_1; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_131 = 6'h2 == L0Index ? io_FromL1 : L0Memory_2; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_132 = 6'h3 == L0Index ? io_FromL1 : L0Memory_3; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_133 = 6'h4 == L0Index ? io_FromL1 : L0Memory_4; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_134 = 6'h5 == L0Index ? io_FromL1 : L0Memory_5; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_135 = 6'h6 == L0Index ? io_FromL1 : L0Memory_6; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_136 = 6'h7 == L0Index ? io_FromL1 : L0Memory_7; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_137 = 6'h8 == L0Index ? io_FromL1 : L0Memory_8; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_138 = 6'h9 == L0Index ? io_FromL1 : L0Memory_9; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_139 = 6'ha == L0Index ? io_FromL1 : L0Memory_10; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_140 = 6'hb == L0Index ? io_FromL1 : L0Memory_11; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_141 = 6'hc == L0Index ? io_FromL1 : L0Memory_12; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_142 = 6'hd == L0Index ? io_FromL1 : L0Memory_13; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_143 = 6'he == L0Index ? io_FromL1 : L0Memory_14; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_144 = 6'hf == L0Index ? io_FromL1 : L0Memory_15; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_145 = 6'h10 == L0Index ? io_FromL1 : L0Memory_16; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_146 = 6'h11 == L0Index ? io_FromL1 : L0Memory_17; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_147 = 6'h12 == L0Index ? io_FromL1 : L0Memory_18; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_148 = 6'h13 == L0Index ? io_FromL1 : L0Memory_19; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_149 = 6'h14 == L0Index ? io_FromL1 : L0Memory_20; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_150 = 6'h15 == L0Index ? io_FromL1 : L0Memory_21; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_151 = 6'h16 == L0Index ? io_FromL1 : L0Memory_22; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_152 = 6'h17 == L0Index ? io_FromL1 : L0Memory_23; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_153 = 6'h18 == L0Index ? io_FromL1 : L0Memory_24; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_154 = 6'h19 == L0Index ? io_FromL1 : L0Memory_25; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_155 = 6'h1a == L0Index ? io_FromL1 : L0Memory_26; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_156 = 6'h1b == L0Index ? io_FromL1 : L0Memory_27; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_157 = 6'h1c == L0Index ? io_FromL1 : L0Memory_28; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_158 = 6'h1d == L0Index ? io_FromL1 : L0Memory_29; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_159 = 6'h1e == L0Index ? io_FromL1 : L0Memory_30; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_160 = 6'h1f == L0Index ? io_FromL1 : L0Memory_31; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_161 = 6'h20 == L0Index ? io_FromL1 : L0Memory_32; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_162 = 6'h21 == L0Index ? io_FromL1 : L0Memory_33; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_163 = 6'h22 == L0Index ? io_FromL1 : L0Memory_34; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_164 = 6'h23 == L0Index ? io_FromL1 : L0Memory_35; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_165 = 6'h24 == L0Index ? io_FromL1 : L0Memory_36; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_166 = 6'h25 == L0Index ? io_FromL1 : L0Memory_37; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_167 = 6'h26 == L0Index ? io_FromL1 : L0Memory_38; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_168 = 6'h27 == L0Index ? io_FromL1 : L0Memory_39; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_169 = 6'h28 == L0Index ? io_FromL1 : L0Memory_40; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_170 = 6'h29 == L0Index ? io_FromL1 : L0Memory_41; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_171 = 6'h2a == L0Index ? io_FromL1 : L0Memory_42; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_172 = 6'h2b == L0Index ? io_FromL1 : L0Memory_43; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_173 = 6'h2c == L0Index ? io_FromL1 : L0Memory_44; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_174 = 6'h2d == L0Index ? io_FromL1 : L0Memory_45; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_175 = 6'h2e == L0Index ? io_FromL1 : L0Memory_46; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_176 = 6'h2f == L0Index ? io_FromL1 : L0Memory_47; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_177 = 6'h30 == L0Index ? io_FromL1 : L0Memory_48; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_178 = 6'h31 == L0Index ? io_FromL1 : L0Memory_49; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_179 = 6'h32 == L0Index ? io_FromL1 : L0Memory_50; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_180 = 6'h33 == L0Index ? io_FromL1 : L0Memory_51; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_181 = 6'h34 == L0Index ? io_FromL1 : L0Memory_52; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_182 = 6'h35 == L0Index ? io_FromL1 : L0Memory_53; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_183 = 6'h36 == L0Index ? io_FromL1 : L0Memory_54; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_184 = 6'h37 == L0Index ? io_FromL1 : L0Memory_55; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_185 = 6'h38 == L0Index ? io_FromL1 : L0Memory_56; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_186 = 6'h39 == L0Index ? io_FromL1 : L0Memory_57; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_187 = 6'h3a == L0Index ? io_FromL1 : L0Memory_58; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_188 = 6'h3b == L0Index ? io_FromL1 : L0Memory_59; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_189 = 6'h3c == L0Index ? io_FromL1 : L0Memory_60; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_190 = 6'h3d == L0Index ? io_FromL1 : L0Memory_61; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_191 = 6'h3e == L0Index ? io_FromL1 : L0Memory_62; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_192 = 6'h3f == L0Index ? io_FromL1 : L0Memory_63; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_193 = 7'h40 == _GEN_793 ? io_FromL1 : L0Memory_64; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_194 = 7'h41 == _GEN_793 ? io_FromL1 : L0Memory_65; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_195 = 7'h42 == _GEN_793 ? io_FromL1 : L0Memory_66; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_196 = 7'h43 == _GEN_793 ? io_FromL1 : L0Memory_67; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_197 = 7'h44 == _GEN_793 ? io_FromL1 : L0Memory_68; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_198 = 7'h45 == _GEN_793 ? io_FromL1 : L0Memory_69; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_199 = 7'h46 == _GEN_793 ? io_FromL1 : L0Memory_70; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_200 = 7'h47 == _GEN_793 ? io_FromL1 : L0Memory_71; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_201 = 7'h48 == _GEN_793 ? io_FromL1 : L0Memory_72; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_202 = 7'h49 == _GEN_793 ? io_FromL1 : L0Memory_73; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_203 = 7'h4a == _GEN_793 ? io_FromL1 : L0Memory_74; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_204 = 7'h4b == _GEN_793 ? io_FromL1 : L0Memory_75; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_205 = 7'h4c == _GEN_793 ? io_FromL1 : L0Memory_76; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_206 = 7'h4d == _GEN_793 ? io_FromL1 : L0Memory_77; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_207 = 7'h4e == _GEN_793 ? io_FromL1 : L0Memory_78; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_208 = 7'h4f == _GEN_793 ? io_FromL1 : L0Memory_79; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_209 = 7'h50 == _GEN_793 ? io_FromL1 : L0Memory_80; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_210 = 7'h51 == _GEN_793 ? io_FromL1 : L0Memory_81; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_211 = 7'h52 == _GEN_793 ? io_FromL1 : L0Memory_82; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_212 = 7'h53 == _GEN_793 ? io_FromL1 : L0Memory_83; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_213 = 7'h54 == _GEN_793 ? io_FromL1 : L0Memory_84; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_214 = 7'h55 == _GEN_793 ? io_FromL1 : L0Memory_85; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_215 = 7'h56 == _GEN_793 ? io_FromL1 : L0Memory_86; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_216 = 7'h57 == _GEN_793 ? io_FromL1 : L0Memory_87; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_217 = 7'h58 == _GEN_793 ? io_FromL1 : L0Memory_88; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_218 = 7'h59 == _GEN_793 ? io_FromL1 : L0Memory_89; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_219 = 7'h5a == _GEN_793 ? io_FromL1 : L0Memory_90; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_220 = 7'h5b == _GEN_793 ? io_FromL1 : L0Memory_91; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_221 = 7'h5c == _GEN_793 ? io_FromL1 : L0Memory_92; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_222 = 7'h5d == _GEN_793 ? io_FromL1 : L0Memory_93; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_223 = 7'h5e == _GEN_793 ? io_FromL1 : L0Memory_94; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_224 = 7'h5f == _GEN_793 ? io_FromL1 : L0Memory_95; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_225 = 7'h60 == _GEN_793 ? io_FromL1 : L0Memory_96; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_226 = 7'h61 == _GEN_793 ? io_FromL1 : L0Memory_97; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_227 = 7'h62 == _GEN_793 ? io_FromL1 : L0Memory_98; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_228 = 7'h63 == _GEN_793 ? io_FromL1 : L0Memory_99; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [5:0] _L0Index_T_2 = L0Index + 6'h1; // @[PEArray.scala 200:28]
  wire [15:0] _GEN_229 = count >= 10'h1 & count <= _T_27 ? _GEN_129 : L0Memory_0; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_230 = count >= 10'h1 & count <= _T_27 ? _GEN_130 : L0Memory_1; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_231 = count >= 10'h1 & count <= _T_27 ? _GEN_131 : L0Memory_2; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_232 = count >= 10'h1 & count <= _T_27 ? _GEN_132 : L0Memory_3; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_233 = count >= 10'h1 & count <= _T_27 ? _GEN_133 : L0Memory_4; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_234 = count >= 10'h1 & count <= _T_27 ? _GEN_134 : L0Memory_5; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_235 = count >= 10'h1 & count <= _T_27 ? _GEN_135 : L0Memory_6; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_236 = count >= 10'h1 & count <= _T_27 ? _GEN_136 : L0Memory_7; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_237 = count >= 10'h1 & count <= _T_27 ? _GEN_137 : L0Memory_8; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_238 = count >= 10'h1 & count <= _T_27 ? _GEN_138 : L0Memory_9; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_239 = count >= 10'h1 & count <= _T_27 ? _GEN_139 : L0Memory_10; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_240 = count >= 10'h1 & count <= _T_27 ? _GEN_140 : L0Memory_11; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_241 = count >= 10'h1 & count <= _T_27 ? _GEN_141 : L0Memory_12; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_242 = count >= 10'h1 & count <= _T_27 ? _GEN_142 : L0Memory_13; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_243 = count >= 10'h1 & count <= _T_27 ? _GEN_143 : L0Memory_14; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_244 = count >= 10'h1 & count <= _T_27 ? _GEN_144 : L0Memory_15; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_245 = count >= 10'h1 & count <= _T_27 ? _GEN_145 : L0Memory_16; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_246 = count >= 10'h1 & count <= _T_27 ? _GEN_146 : L0Memory_17; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_247 = count >= 10'h1 & count <= _T_27 ? _GEN_147 : L0Memory_18; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_248 = count >= 10'h1 & count <= _T_27 ? _GEN_148 : L0Memory_19; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_249 = count >= 10'h1 & count <= _T_27 ? _GEN_149 : L0Memory_20; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_250 = count >= 10'h1 & count <= _T_27 ? _GEN_150 : L0Memory_21; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_251 = count >= 10'h1 & count <= _T_27 ? _GEN_151 : L0Memory_22; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_252 = count >= 10'h1 & count <= _T_27 ? _GEN_152 : L0Memory_23; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_253 = count >= 10'h1 & count <= _T_27 ? _GEN_153 : L0Memory_24; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_254 = count >= 10'h1 & count <= _T_27 ? _GEN_154 : L0Memory_25; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_255 = count >= 10'h1 & count <= _T_27 ? _GEN_155 : L0Memory_26; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_256 = count >= 10'h1 & count <= _T_27 ? _GEN_156 : L0Memory_27; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_257 = count >= 10'h1 & count <= _T_27 ? _GEN_157 : L0Memory_28; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_258 = count >= 10'h1 & count <= _T_27 ? _GEN_158 : L0Memory_29; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_259 = count >= 10'h1 & count <= _T_27 ? _GEN_159 : L0Memory_30; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_260 = count >= 10'h1 & count <= _T_27 ? _GEN_160 : L0Memory_31; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_261 = count >= 10'h1 & count <= _T_27 ? _GEN_161 : L0Memory_32; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_262 = count >= 10'h1 & count <= _T_27 ? _GEN_162 : L0Memory_33; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_263 = count >= 10'h1 & count <= _T_27 ? _GEN_163 : L0Memory_34; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_264 = count >= 10'h1 & count <= _T_27 ? _GEN_164 : L0Memory_35; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_265 = count >= 10'h1 & count <= _T_27 ? _GEN_165 : L0Memory_36; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_266 = count >= 10'h1 & count <= _T_27 ? _GEN_166 : L0Memory_37; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_267 = count >= 10'h1 & count <= _T_27 ? _GEN_167 : L0Memory_38; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_268 = count >= 10'h1 & count <= _T_27 ? _GEN_168 : L0Memory_39; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_269 = count >= 10'h1 & count <= _T_27 ? _GEN_169 : L0Memory_40; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_270 = count >= 10'h1 & count <= _T_27 ? _GEN_170 : L0Memory_41; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_271 = count >= 10'h1 & count <= _T_27 ? _GEN_171 : L0Memory_42; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_272 = count >= 10'h1 & count <= _T_27 ? _GEN_172 : L0Memory_43; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_273 = count >= 10'h1 & count <= _T_27 ? _GEN_173 : L0Memory_44; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_274 = count >= 10'h1 & count <= _T_27 ? _GEN_174 : L0Memory_45; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_275 = count >= 10'h1 & count <= _T_27 ? _GEN_175 : L0Memory_46; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_276 = count >= 10'h1 & count <= _T_27 ? _GEN_176 : L0Memory_47; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_277 = count >= 10'h1 & count <= _T_27 ? _GEN_177 : L0Memory_48; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_278 = count >= 10'h1 & count <= _T_27 ? _GEN_178 : L0Memory_49; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_279 = count >= 10'h1 & count <= _T_27 ? _GEN_179 : L0Memory_50; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_280 = count >= 10'h1 & count <= _T_27 ? _GEN_180 : L0Memory_51; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_281 = count >= 10'h1 & count <= _T_27 ? _GEN_181 : L0Memory_52; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_282 = count >= 10'h1 & count <= _T_27 ? _GEN_182 : L0Memory_53; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_283 = count >= 10'h1 & count <= _T_27 ? _GEN_183 : L0Memory_54; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_284 = count >= 10'h1 & count <= _T_27 ? _GEN_184 : L0Memory_55; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_285 = count >= 10'h1 & count <= _T_27 ? _GEN_185 : L0Memory_56; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_286 = count >= 10'h1 & count <= _T_27 ? _GEN_186 : L0Memory_57; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_287 = count >= 10'h1 & count <= _T_27 ? _GEN_187 : L0Memory_58; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_288 = count >= 10'h1 & count <= _T_27 ? _GEN_188 : L0Memory_59; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_289 = count >= 10'h1 & count <= _T_27 ? _GEN_189 : L0Memory_60; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_290 = count >= 10'h1 & count <= _T_27 ? _GEN_190 : L0Memory_61; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_291 = count >= 10'h1 & count <= _T_27 ? _GEN_191 : L0Memory_62; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_292 = count >= 10'h1 & count <= _T_27 ? _GEN_192 : L0Memory_63; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_293 = count >= 10'h1 & count <= _T_27 ? _GEN_193 : L0Memory_64; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_294 = count >= 10'h1 & count <= _T_27 ? _GEN_194 : L0Memory_65; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_295 = count >= 10'h1 & count <= _T_27 ? _GEN_195 : L0Memory_66; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_296 = count >= 10'h1 & count <= _T_27 ? _GEN_196 : L0Memory_67; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_297 = count >= 10'h1 & count <= _T_27 ? _GEN_197 : L0Memory_68; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_298 = count >= 10'h1 & count <= _T_27 ? _GEN_198 : L0Memory_69; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_299 = count >= 10'h1 & count <= _T_27 ? _GEN_199 : L0Memory_70; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_300 = count >= 10'h1 & count <= _T_27 ? _GEN_200 : L0Memory_71; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_301 = count >= 10'h1 & count <= _T_27 ? _GEN_201 : L0Memory_72; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_302 = count >= 10'h1 & count <= _T_27 ? _GEN_202 : L0Memory_73; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_303 = count >= 10'h1 & count <= _T_27 ? _GEN_203 : L0Memory_74; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_304 = count >= 10'h1 & count <= _T_27 ? _GEN_204 : L0Memory_75; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_305 = count >= 10'h1 & count <= _T_27 ? _GEN_205 : L0Memory_76; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_306 = count >= 10'h1 & count <= _T_27 ? _GEN_206 : L0Memory_77; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_307 = count >= 10'h1 & count <= _T_27 ? _GEN_207 : L0Memory_78; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_308 = count >= 10'h1 & count <= _T_27 ? _GEN_208 : L0Memory_79; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_309 = count >= 10'h1 & count <= _T_27 ? _GEN_209 : L0Memory_80; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_310 = count >= 10'h1 & count <= _T_27 ? _GEN_210 : L0Memory_81; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_311 = count >= 10'h1 & count <= _T_27 ? _GEN_211 : L0Memory_82; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_312 = count >= 10'h1 & count <= _T_27 ? _GEN_212 : L0Memory_83; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_313 = count >= 10'h1 & count <= _T_27 ? _GEN_213 : L0Memory_84; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_314 = count >= 10'h1 & count <= _T_27 ? _GEN_214 : L0Memory_85; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_315 = count >= 10'h1 & count <= _T_27 ? _GEN_215 : L0Memory_86; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_316 = count >= 10'h1 & count <= _T_27 ? _GEN_216 : L0Memory_87; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_317 = count >= 10'h1 & count <= _T_27 ? _GEN_217 : L0Memory_88; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_318 = count >= 10'h1 & count <= _T_27 ? _GEN_218 : L0Memory_89; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_319 = count >= 10'h1 & count <= _T_27 ? _GEN_219 : L0Memory_90; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_320 = count >= 10'h1 & count <= _T_27 ? _GEN_220 : L0Memory_91; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_321 = count >= 10'h1 & count <= _T_27 ? _GEN_221 : L0Memory_92; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_322 = count >= 10'h1 & count <= _T_27 ? _GEN_222 : L0Memory_93; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_323 = count >= 10'h1 & count <= _T_27 ? _GEN_223 : L0Memory_94; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_324 = count >= 10'h1 & count <= _T_27 ? _GEN_224 : L0Memory_95; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_325 = count >= 10'h1 & count <= _T_27 ? _GEN_225 : L0Memory_96; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_326 = count >= 10'h1 & count <= _T_27 ? _GEN_226 : L0Memory_97; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_327 = count >= 10'h1 & count <= _T_27 ? _GEN_227 : L0Memory_98; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_328 = count >= 10'h1 & count <= _T_27 ? _GEN_228 : L0Memory_99; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [5:0] _GEN_329 = count >= 10'h1 & count <= _T_27 ? _L0Index_T_2 : _GEN_128; // @[PEArray.scala 198:59 PEArray.scala 200:17]
  wire [9:0] _GEN_330 = count == count_max ? 10'h0 : _GEN_127; // @[PEArray.scala 202:32 PEArray.scala 203:15]
  wire [2:0] _GEN_331 = count == count_max ? 3'h0 : state; // @[PEArray.scala 202:32 PEArray.scala 204:15 PEArray.scala 100:22]
  wire [9:0] _GEN_865 = {{4'd0}, GRU_out_width}; // @[PEArray.scala 220:19]
  wire [9:0] _GEN_0 = count % _GEN_865; // @[PEArray.scala 220:19]
  wire [5:0] _T_36 = _GEN_0[5:0]; // @[PEArray.scala 220:19]
  wire [5:0] _T_38 = GRU_out_width - 6'h1; // @[PEArray.scala 220:55]
  wire [5:0] _GEN_334 = _T_36 == _T_38 ? _L0Index_T_2 : L0index_begin; // @[PEArray.scala 220:62 PEArray.scala 221:17 PEArray.scala 214:15]
  wire [5:0] _GEN_346 = _T_41 ? _GEN_334 : L0Index; // @[Conditional.scala 39:67 PEArray.scala 39:24]
  wire [9:0] _GEN_347 = _T_41 ? _GEN_330 : count; // @[Conditional.scala 39:67 PEArray.scala 101:22]
  wire [2:0] _GEN_348 = _T_41 ? _GEN_331 : state; // @[Conditional.scala 39:67 PEArray.scala 100:22]
  wire [5:0] _GEN_353 = _T_31 ? _GEN_334 : _GEN_346; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_354 = _T_31 ? _GEN_330 : _GEN_347; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_355 = _T_31 ? _GEN_331 : _GEN_348; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_356 = _T_22 ? _GEN_330 : _GEN_354; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_357 = _T_22 ? _GEN_329 : _GEN_353; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_458 = _T_22 ? _GEN_331 : _GEN_355; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_690 = _T_3 ? _GEN_118 : {{2'd0}, GRU_out_width}; // @[Conditional.scala 40:58 PEArray.scala 104:26]
  FP16MulAdder FP16MAC ( // @[PEArray.scala 72:23]
    .io_a(FP16MAC_io_a),
    .io_b(FP16MAC_io_b),
    .io_c(FP16MAC_io_c),
    .io_out(FP16MAC_io_out)
  );
  assign io_ToRightPE = mux3out_reg; // @[PEArray.scala 95:16]
  assign io_ToBelowPE = mux2out_reg; // @[PEArray.scala 94:16]
  assign FP16MAC_io_a = sel1 ? io_FromL1 : io_FromLeftPE; // @[PEArray.scala 50:14 PEArray.scala 50:23 PEArray.scala 51:24]
  assign FP16MAC_io_b = sel5 ? mux4out : _GEN_105; // @[PEArray.scala 77:13 PEArray.scala 78:18 PEArray.scala 81:18]
  assign FP16MAC_io_c = sel5 ? _GEN_105 : mux4out; // @[PEArray.scala 77:13 PEArray.scala 79:18 PEArray.scala 82:18]
  always @(posedge clock) begin
    if (reset) begin // @[PEArray.scala 39:24]
      L0Index <= 6'h0; // @[PEArray.scala 39:24]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h2; // @[PEArray.scala 159:15]
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        L0Index <= 6'hd; // @[PEArray.scala 181:15]
      end else begin
        L0Index <= _GEN_357;
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_0 <= _GEN_229;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_1 <= _GEN_230;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_2 <= _GEN_231;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_3 <= _GEN_232;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_4 <= _GEN_233;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_5 <= _GEN_234;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_6 <= _GEN_235;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_7 <= _GEN_236;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_8 <= _GEN_237;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_9 <= _GEN_238;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_10 <= _GEN_239;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_11 <= _GEN_240;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_12 <= _GEN_241;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_13 <= _GEN_242;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_14 <= _GEN_243;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_15 <= _GEN_244;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_16 <= _GEN_245;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_17 <= _GEN_246;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_18 <= _GEN_247;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_19 <= _GEN_248;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_20 <= _GEN_249;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_21 <= _GEN_250;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_22 <= _GEN_251;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_23 <= _GEN_252;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_24 <= _GEN_253;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_25 <= _GEN_254;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_26 <= _GEN_255;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_27 <= _GEN_256;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_28 <= _GEN_257;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_29 <= _GEN_258;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_30 <= _GEN_259;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_31 <= _GEN_260;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_32 <= _GEN_261;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_33 <= _GEN_262;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_34 <= _GEN_263;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_35 <= _GEN_264;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_36 <= _GEN_265;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_37 <= _GEN_266;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_38 <= _GEN_267;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_39 <= _GEN_268;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_40 <= _GEN_269;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_41 <= _GEN_270;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_42 <= _GEN_271;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_43 <= _GEN_272;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_44 <= _GEN_273;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_45 <= _GEN_274;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_46 <= _GEN_275;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_47 <= _GEN_276;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_48 <= _GEN_277;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_49 <= _GEN_278;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_50 <= _GEN_279;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_51 <= _GEN_280;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_52 <= _GEN_281;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_53 <= _GEN_282;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_54 <= _GEN_283;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_55 <= _GEN_284;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_56 <= _GEN_285;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_57 <= _GEN_286;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_58 <= _GEN_287;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_59 <= _GEN_288;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_60 <= _GEN_289;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_61 <= _GEN_290;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_62 <= _GEN_291;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_63 <= _GEN_292;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_64 <= _GEN_293;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_65 <= _GEN_294;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_66 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_67 <= _GEN_296;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_68 <= _GEN_297;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_69 <= _GEN_298;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_70 <= _GEN_299;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_71 <= _GEN_300;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_72 <= _GEN_301;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_73 <= _GEN_302;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_74 <= _GEN_303;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_75 <= _GEN_304;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_76 <= _GEN_305;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_77 <= _GEN_306;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_78 <= _GEN_307;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_79 <= _GEN_308;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_80 <= _GEN_309;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_81 <= _GEN_310;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_82 <= _GEN_311;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_83 <= _GEN_312;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_84 <= _GEN_313;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_85 <= _GEN_314;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_86 <= _GEN_315;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_87 <= _GEN_316;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_88 <= _GEN_317;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_89 <= _GEN_318;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_90 <= _GEN_319;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_91 <= _GEN_320;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_92 <= _GEN_321;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_93 <= _GEN_322;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_94 <= _GEN_323;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_95 <= _GEN_324;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_96 <= _GEN_325;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_97 <= _GEN_326;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_98 <= _GEN_327;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_99 <= _GEN_328;
          end
        end
      end
    end
    if (reset) begin // @[PEArray.scala 100:22]
      state <= 3'h0; // @[PEArray.scala 100:22]
    end else if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[1]) begin // @[PEArray.scala 116:57]
        if (_T_6) begin // @[Conditional.scala 40:58]
          state <= 3'h0; // @[PEArray.scala 120:19]
        end else begin
          state <= _GEN_113;
        end
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      if (count == 10'h33) begin // @[PEArray.scala 164:27]
        state <= 3'h0; // @[PEArray.scala 166:15]
      end
    end else if (_T_16) begin // @[Conditional.scala 39:67]
      state <= _GEN_126;
    end else begin
      state <= _GEN_458;
    end
    if (reset) begin // @[PEArray.scala 90:28]
      mux2out_reg <= 16'h0; // @[PEArray.scala 90:28]
    end else begin
      mux2out_reg <= MAC_out; // @[PEArray.scala 90:28]
    end
    if (reset) begin // @[PEArray.scala 91:28]
      mux3out_reg <= 16'h0; // @[PEArray.scala 91:28]
    end else if (sel3) begin // @[PEArray.scala 56:14]
      mux3out_reg <= MAC_out; // @[PEArray.scala 56:23]
    end else if (sel1) begin // @[PEArray.scala 50:14]
      mux3out_reg <= io_FromL1; // @[PEArray.scala 50:23]
    end else begin
      mux3out_reg <= io_FromLeftPE; // @[PEArray.scala 51:24]
    end
    if (reset) begin // @[PEArray.scala 101:22]
      count <= 10'h0; // @[PEArray.scala 101:22]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        if (count == 10'h33) begin // @[PEArray.scala 164:27]
          count <= 10'h0; // @[PEArray.scala 165:15]
        end else begin
          count <= _GEN_120;
        end
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        count <= _GEN_125;
      end else begin
        count <= _GEN_356;
      end
    end
    if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[1]) begin // @[PEArray.scala 116:57]
        count_max <= io_control_signal_count; // @[PEArray.scala 143:19]
      end
    end
    if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[1]) begin // @[PEArray.scala 116:57]
        L0index_begin <= io_control_signal_L0index; // @[PEArray.scala 144:23]
      end
    end
    GRU_out_width <= _GEN_690[5:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  L0Index = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  L0Memory_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  L0Memory_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  L0Memory_2 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  L0Memory_3 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  L0Memory_4 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  L0Memory_5 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  L0Memory_6 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  L0Memory_7 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  L0Memory_8 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  L0Memory_9 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  L0Memory_10 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  L0Memory_11 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  L0Memory_12 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  L0Memory_13 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  L0Memory_14 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  L0Memory_15 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  L0Memory_16 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  L0Memory_17 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  L0Memory_18 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  L0Memory_19 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  L0Memory_20 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  L0Memory_21 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  L0Memory_22 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  L0Memory_23 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  L0Memory_24 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  L0Memory_25 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  L0Memory_26 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  L0Memory_27 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  L0Memory_28 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  L0Memory_29 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  L0Memory_30 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  L0Memory_31 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  L0Memory_32 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  L0Memory_33 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  L0Memory_34 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  L0Memory_35 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  L0Memory_36 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  L0Memory_37 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  L0Memory_38 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  L0Memory_39 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  L0Memory_40 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  L0Memory_41 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  L0Memory_42 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  L0Memory_43 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  L0Memory_44 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  L0Memory_45 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  L0Memory_46 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  L0Memory_47 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  L0Memory_48 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  L0Memory_49 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  L0Memory_50 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  L0Memory_51 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  L0Memory_52 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  L0Memory_53 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  L0Memory_54 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  L0Memory_55 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  L0Memory_56 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  L0Memory_57 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  L0Memory_58 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  L0Memory_59 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  L0Memory_60 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  L0Memory_61 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  L0Memory_62 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  L0Memory_63 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  L0Memory_64 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  L0Memory_65 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  L0Memory_66 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  L0Memory_67 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  L0Memory_68 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  L0Memory_69 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  L0Memory_70 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  L0Memory_71 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  L0Memory_72 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  L0Memory_73 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  L0Memory_74 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  L0Memory_75 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  L0Memory_76 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  L0Memory_77 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  L0Memory_78 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  L0Memory_79 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  L0Memory_80 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  L0Memory_81 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  L0Memory_82 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  L0Memory_83 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  L0Memory_84 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  L0Memory_85 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  L0Memory_86 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  L0Memory_87 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  L0Memory_88 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  L0Memory_89 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  L0Memory_90 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  L0Memory_91 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  L0Memory_92 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  L0Memory_93 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  L0Memory_94 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  L0Memory_95 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  L0Memory_96 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  L0Memory_97 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  L0Memory_98 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  L0Memory_99 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  state = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  mux2out_reg = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  mux3out_reg = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  count = _RAND_104[9:0];
  _RAND_105 = {1{`RANDOM}};
  count_max = _RAND_105[9:0];
  _RAND_106 = {1{`RANDOM}};
  L0index_begin = _RAND_106[5:0];
  _RAND_107 = {1{`RANDOM}};
  GRU_out_width = _RAND_107[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PE_33(
  input         clock,
  input         reset,
  input  [15:0] io_FromAbovePE,
  input  [15:0] io_FromLeftPE,
  input  [15:0] io_FromL1,
  input  [11:0] io_control_signal_mask,
  output [15:0] io_ToBelowPE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] FP16MAC_io_a; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_b; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_c; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_out; // @[PEArray.scala 72:23]
  reg [5:0] L0Index; // @[PEArray.scala 39:24]
  reg [15:0] L0Memory_0; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_1; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_2; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_3; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_4; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_5; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_6; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_7; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_8; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_9; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_10; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_11; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_12; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_13; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_14; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_15; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_16; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_17; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_18; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_19; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_20; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_21; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_22; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_23; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_24; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_25; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_26; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_27; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_28; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_29; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_30; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_31; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_32; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_33; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_34; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_35; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_36; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_37; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_38; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_39; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_40; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_41; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_42; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_43; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_44; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_45; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_46; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_47; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_48; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_49; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_50; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_51; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_52; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_53; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_54; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_55; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_56; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_57; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_58; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_59; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_60; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_61; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_62; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_63; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_64; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_65; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_66; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_67; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_68; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_69; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_70; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_71; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_72; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_73; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_74; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_75; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_76; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_77; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_78; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_79; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_80; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_81; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_82; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_83; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_84; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_85; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_86; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_87; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_88; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_89; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_90; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_91; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_92; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_93; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_94; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_95; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_96; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_97; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_98; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_99; // @[PEArray.scala 40:21]
  reg [2:0] state; // @[PEArray.scala 100:22]
  wire  _T_3 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_12 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_16 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_22 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_31 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_41 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_342 = _T_41 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 231:12 PEArray.scala 32:8]
  wire  _GEN_349 = _T_31 ? 1'h0 : _GEN_342; // @[Conditional.scala 39:67 PEArray.scala 208:12]
  wire  _GEN_459 = _T_22 | _GEN_349; // @[Conditional.scala 39:67 PEArray.scala 32:8]
  wire  _GEN_463 = _T_16 ? 1'h0 : _GEN_459; // @[Conditional.scala 39:67]
  wire  _GEN_572 = _T_12 | _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 149:12]
  wire  sel1 = _T_3 | _GEN_572; // @[Conditional.scala 40:58 PEArray.scala 108:12]
  wire [15:0] MAC_out = FP16MAC_io_out; // @[PEArray.scala 47:21 PEArray.scala 85:11]
  wire [1:0] _GEN_344 = _T_41 ? 2'h2 : 2'h0; // @[Conditional.scala 39:67 PEArray.scala 233:12 PEArray.scala 35:8]
  wire [1:0] _GEN_351 = _T_31 ? 2'h2 : _GEN_344; // @[Conditional.scala 39:67 PEArray.scala 210:12]
  wire [1:0] _GEN_461 = _T_22 ? 2'h0 : _GEN_351; // @[Conditional.scala 39:67 PEArray.scala 35:8]
  wire [1:0] _GEN_466 = _T_16 ? 2'h0 : _GEN_461; // @[Conditional.scala 39:67 PEArray.scala 178:12]
  wire [1:0] _GEN_574 = _T_12 ? 2'h0 : _GEN_466; // @[Conditional.scala 39:67]
  wire [1:0] sel4 = _T_3 ? 2'h0 : _GEN_574; // @[Conditional.scala 40:58 PEArray.scala 111:12]
  wire [15:0] _GEN_3 = sel4 == 2'h2 ? io_FromL1 : 16'h0; // @[PEArray.scala 65:28 PEArray.scala 66:15 PEArray.scala 69:15]
  wire [15:0] _GEN_4 = sel4 == 2'h1 ? io_FromAbovePE : _GEN_3; // @[PEArray.scala 62:28 PEArray.scala 63:15]
  wire [15:0] mux4out = sel4 == 2'h0 ? 16'h0 : _GEN_4; // @[PEArray.scala 59:22 PEArray.scala 60:13]
  wire [15:0] _GEN_7 = 6'h1 == L0Index ? L0Memory_1 : L0Memory_0; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_8 = 6'h2 == L0Index ? L0Memory_2 : _GEN_7; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_9 = 6'h3 == L0Index ? L0Memory_3 : _GEN_8; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_10 = 6'h4 == L0Index ? L0Memory_4 : _GEN_9; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_11 = 6'h5 == L0Index ? L0Memory_5 : _GEN_10; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_12 = 6'h6 == L0Index ? L0Memory_6 : _GEN_11; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_13 = 6'h7 == L0Index ? L0Memory_7 : _GEN_12; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_14 = 6'h8 == L0Index ? L0Memory_8 : _GEN_13; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_15 = 6'h9 == L0Index ? L0Memory_9 : _GEN_14; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_16 = 6'ha == L0Index ? L0Memory_10 : _GEN_15; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_17 = 6'hb == L0Index ? L0Memory_11 : _GEN_16; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_18 = 6'hc == L0Index ? L0Memory_12 : _GEN_17; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_19 = 6'hd == L0Index ? L0Memory_13 : _GEN_18; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_20 = 6'he == L0Index ? L0Memory_14 : _GEN_19; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_21 = 6'hf == L0Index ? L0Memory_15 : _GEN_20; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_22 = 6'h10 == L0Index ? L0Memory_16 : _GEN_21; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_23 = 6'h11 == L0Index ? L0Memory_17 : _GEN_22; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_24 = 6'h12 == L0Index ? L0Memory_18 : _GEN_23; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_25 = 6'h13 == L0Index ? L0Memory_19 : _GEN_24; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_26 = 6'h14 == L0Index ? L0Memory_20 : _GEN_25; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_27 = 6'h15 == L0Index ? L0Memory_21 : _GEN_26; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_28 = 6'h16 == L0Index ? L0Memory_22 : _GEN_27; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_29 = 6'h17 == L0Index ? L0Memory_23 : _GEN_28; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_30 = 6'h18 == L0Index ? L0Memory_24 : _GEN_29; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_31 = 6'h19 == L0Index ? L0Memory_25 : _GEN_30; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_32 = 6'h1a == L0Index ? L0Memory_26 : _GEN_31; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_33 = 6'h1b == L0Index ? L0Memory_27 : _GEN_32; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_34 = 6'h1c == L0Index ? L0Memory_28 : _GEN_33; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_35 = 6'h1d == L0Index ? L0Memory_29 : _GEN_34; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_36 = 6'h1e == L0Index ? L0Memory_30 : _GEN_35; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_37 = 6'h1f == L0Index ? L0Memory_31 : _GEN_36; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_38 = 6'h20 == L0Index ? L0Memory_32 : _GEN_37; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_39 = 6'h21 == L0Index ? L0Memory_33 : _GEN_38; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_40 = 6'h22 == L0Index ? L0Memory_34 : _GEN_39; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_41 = 6'h23 == L0Index ? L0Memory_35 : _GEN_40; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_42 = 6'h24 == L0Index ? L0Memory_36 : _GEN_41; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_43 = 6'h25 == L0Index ? L0Memory_37 : _GEN_42; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_44 = 6'h26 == L0Index ? L0Memory_38 : _GEN_43; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_45 = 6'h27 == L0Index ? L0Memory_39 : _GEN_44; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_46 = 6'h28 == L0Index ? L0Memory_40 : _GEN_45; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_47 = 6'h29 == L0Index ? L0Memory_41 : _GEN_46; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_48 = 6'h2a == L0Index ? L0Memory_42 : _GEN_47; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_49 = 6'h2b == L0Index ? L0Memory_43 : _GEN_48; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_50 = 6'h2c == L0Index ? L0Memory_44 : _GEN_49; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_51 = 6'h2d == L0Index ? L0Memory_45 : _GEN_50; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_52 = 6'h2e == L0Index ? L0Memory_46 : _GEN_51; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_53 = 6'h2f == L0Index ? L0Memory_47 : _GEN_52; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_54 = 6'h30 == L0Index ? L0Memory_48 : _GEN_53; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_55 = 6'h31 == L0Index ? L0Memory_49 : _GEN_54; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_56 = 6'h32 == L0Index ? L0Memory_50 : _GEN_55; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_57 = 6'h33 == L0Index ? L0Memory_51 : _GEN_56; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_58 = 6'h34 == L0Index ? L0Memory_52 : _GEN_57; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_59 = 6'h35 == L0Index ? L0Memory_53 : _GEN_58; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_60 = 6'h36 == L0Index ? L0Memory_54 : _GEN_59; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_61 = 6'h37 == L0Index ? L0Memory_55 : _GEN_60; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_62 = 6'h38 == L0Index ? L0Memory_56 : _GEN_61; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_63 = 6'h39 == L0Index ? L0Memory_57 : _GEN_62; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_64 = 6'h3a == L0Index ? L0Memory_58 : _GEN_63; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_65 = 6'h3b == L0Index ? L0Memory_59 : _GEN_64; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_66 = 6'h3c == L0Index ? L0Memory_60 : _GEN_65; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_67 = 6'h3d == L0Index ? L0Memory_61 : _GEN_66; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_68 = 6'h3e == L0Index ? L0Memory_62 : _GEN_67; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_69 = 6'h3f == L0Index ? L0Memory_63 : _GEN_68; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [6:0] _GEN_793 = {{1'd0}, L0Index}; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_70 = 7'h40 == _GEN_793 ? L0Memory_64 : _GEN_69; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_71 = 7'h41 == _GEN_793 ? L0Memory_65 : _GEN_70; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_72 = 7'h42 == _GEN_793 ? L0Memory_66 : _GEN_71; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_73 = 7'h43 == _GEN_793 ? L0Memory_67 : _GEN_72; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_74 = 7'h44 == _GEN_793 ? L0Memory_68 : _GEN_73; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_75 = 7'h45 == _GEN_793 ? L0Memory_69 : _GEN_74; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_76 = 7'h46 == _GEN_793 ? L0Memory_70 : _GEN_75; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_77 = 7'h47 == _GEN_793 ? L0Memory_71 : _GEN_76; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_78 = 7'h48 == _GEN_793 ? L0Memory_72 : _GEN_77; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_79 = 7'h49 == _GEN_793 ? L0Memory_73 : _GEN_78; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_80 = 7'h4a == _GEN_793 ? L0Memory_74 : _GEN_79; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_81 = 7'h4b == _GEN_793 ? L0Memory_75 : _GEN_80; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_82 = 7'h4c == _GEN_793 ? L0Memory_76 : _GEN_81; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_83 = 7'h4d == _GEN_793 ? L0Memory_77 : _GEN_82; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_84 = 7'h4e == _GEN_793 ? L0Memory_78 : _GEN_83; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_85 = 7'h4f == _GEN_793 ? L0Memory_79 : _GEN_84; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_86 = 7'h50 == _GEN_793 ? L0Memory_80 : _GEN_85; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_87 = 7'h51 == _GEN_793 ? L0Memory_81 : _GEN_86; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_88 = 7'h52 == _GEN_793 ? L0Memory_82 : _GEN_87; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_89 = 7'h53 == _GEN_793 ? L0Memory_83 : _GEN_88; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_90 = 7'h54 == _GEN_793 ? L0Memory_84 : _GEN_89; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_91 = 7'h55 == _GEN_793 ? L0Memory_85 : _GEN_90; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_92 = 7'h56 == _GEN_793 ? L0Memory_86 : _GEN_91; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_93 = 7'h57 == _GEN_793 ? L0Memory_87 : _GEN_92; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_94 = 7'h58 == _GEN_793 ? L0Memory_88 : _GEN_93; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_95 = 7'h59 == _GEN_793 ? L0Memory_89 : _GEN_94; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_96 = 7'h5a == _GEN_793 ? L0Memory_90 : _GEN_95; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_97 = 7'h5b == _GEN_793 ? L0Memory_91 : _GEN_96; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_98 = 7'h5c == _GEN_793 ? L0Memory_92 : _GEN_97; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_99 = 7'h5d == _GEN_793 ? L0Memory_93 : _GEN_98; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_100 = 7'h5e == _GEN_793 ? L0Memory_94 : _GEN_99; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_101 = 7'h5f == _GEN_793 ? L0Memory_95 : _GEN_100; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_102 = 7'h60 == _GEN_793 ? L0Memory_96 : _GEN_101; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_103 = 7'h61 == _GEN_793 ? L0Memory_97 : _GEN_102; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_104 = 7'h62 == _GEN_793 ? L0Memory_98 : _GEN_103; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_105 = 7'h63 == _GEN_793 ? L0Memory_99 : _GEN_104; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire  _GEN_575 = _T_12 ? 1'h0 : _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 157:12]
  wire  sel5 = _T_3 ? 1'h0 : _GEN_575; // @[Conditional.scala 40:58 PEArray.scala 112:12]
  reg [15:0] mux2out_reg; // @[PEArray.scala 90:28]
  reg [9:0] count; // @[PEArray.scala 101:22]
  reg [5:0] GRU_out_width; // @[PEArray.scala 104:26]
  wire [7:0] _GEN_118 = io_control_signal_mask[0] ? 8'h0 : {{2'd0}, GRU_out_width}; // @[PEArray.scala 116:57 PEArray.scala 145:23 PEArray.scala 104:26]
  wire [9:0] _count_T_1 = count + 10'h1; // @[PEArray.scala 162:24]
  wire [9:0] _GEN_120 = count != 10'h33 ? _count_T_1 : count; // @[PEArray.scala 161:27 PEArray.scala 162:15 PEArray.scala 101:22]
  wire [9:0] _GEN_124 = count != 10'h188 ? _count_T_1 : count; // @[PEArray.scala 183:28 PEArray.scala 184:15 PEArray.scala 101:22]
  wire [9:0] _GEN_125 = count == 10'h188 ? 10'h0 : _GEN_124; // @[PEArray.scala 186:28 PEArray.scala 187:15]
  wire [2:0] _GEN_126 = count == 10'h188 ? 3'h0 : state; // @[PEArray.scala 186:28 PEArray.scala 188:15 PEArray.scala 100:22]
  wire [9:0] _GEN_127 = count != 10'h0 ? _count_T_1 : count; // @[PEArray.scala 192:32 PEArray.scala 193:15 PEArray.scala 101:22]
  wire  _T_24 = count == 10'h0; // @[PEArray.scala 195:18]
  wire [5:0] _GEN_128 = count == 10'h0 ? 6'h0 : L0Index; // @[PEArray.scala 195:26 PEArray.scala 196:17 PEArray.scala 39:24]
  wire [9:0] _T_27 = 10'h0 - 10'h1; // @[PEArray.scala 198:51]
  wire [15:0] _GEN_129 = 6'h0 == L0Index ? io_FromL1 : L0Memory_0; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_130 = 6'h1 == L0Index ? io_FromL1 : L0Memory_1; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_131 = 6'h2 == L0Index ? io_FromL1 : L0Memory_2; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_132 = 6'h3 == L0Index ? io_FromL1 : L0Memory_3; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_133 = 6'h4 == L0Index ? io_FromL1 : L0Memory_4; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_134 = 6'h5 == L0Index ? io_FromL1 : L0Memory_5; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_135 = 6'h6 == L0Index ? io_FromL1 : L0Memory_6; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_136 = 6'h7 == L0Index ? io_FromL1 : L0Memory_7; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_137 = 6'h8 == L0Index ? io_FromL1 : L0Memory_8; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_138 = 6'h9 == L0Index ? io_FromL1 : L0Memory_9; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_139 = 6'ha == L0Index ? io_FromL1 : L0Memory_10; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_140 = 6'hb == L0Index ? io_FromL1 : L0Memory_11; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_141 = 6'hc == L0Index ? io_FromL1 : L0Memory_12; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_142 = 6'hd == L0Index ? io_FromL1 : L0Memory_13; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_143 = 6'he == L0Index ? io_FromL1 : L0Memory_14; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_144 = 6'hf == L0Index ? io_FromL1 : L0Memory_15; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_145 = 6'h10 == L0Index ? io_FromL1 : L0Memory_16; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_146 = 6'h11 == L0Index ? io_FromL1 : L0Memory_17; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_147 = 6'h12 == L0Index ? io_FromL1 : L0Memory_18; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_148 = 6'h13 == L0Index ? io_FromL1 : L0Memory_19; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_149 = 6'h14 == L0Index ? io_FromL1 : L0Memory_20; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_150 = 6'h15 == L0Index ? io_FromL1 : L0Memory_21; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_151 = 6'h16 == L0Index ? io_FromL1 : L0Memory_22; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_152 = 6'h17 == L0Index ? io_FromL1 : L0Memory_23; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_153 = 6'h18 == L0Index ? io_FromL1 : L0Memory_24; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_154 = 6'h19 == L0Index ? io_FromL1 : L0Memory_25; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_155 = 6'h1a == L0Index ? io_FromL1 : L0Memory_26; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_156 = 6'h1b == L0Index ? io_FromL1 : L0Memory_27; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_157 = 6'h1c == L0Index ? io_FromL1 : L0Memory_28; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_158 = 6'h1d == L0Index ? io_FromL1 : L0Memory_29; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_159 = 6'h1e == L0Index ? io_FromL1 : L0Memory_30; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_160 = 6'h1f == L0Index ? io_FromL1 : L0Memory_31; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_161 = 6'h20 == L0Index ? io_FromL1 : L0Memory_32; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_162 = 6'h21 == L0Index ? io_FromL1 : L0Memory_33; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_163 = 6'h22 == L0Index ? io_FromL1 : L0Memory_34; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_164 = 6'h23 == L0Index ? io_FromL1 : L0Memory_35; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_165 = 6'h24 == L0Index ? io_FromL1 : L0Memory_36; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_166 = 6'h25 == L0Index ? io_FromL1 : L0Memory_37; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_167 = 6'h26 == L0Index ? io_FromL1 : L0Memory_38; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_168 = 6'h27 == L0Index ? io_FromL1 : L0Memory_39; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_169 = 6'h28 == L0Index ? io_FromL1 : L0Memory_40; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_170 = 6'h29 == L0Index ? io_FromL1 : L0Memory_41; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_171 = 6'h2a == L0Index ? io_FromL1 : L0Memory_42; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_172 = 6'h2b == L0Index ? io_FromL1 : L0Memory_43; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_173 = 6'h2c == L0Index ? io_FromL1 : L0Memory_44; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_174 = 6'h2d == L0Index ? io_FromL1 : L0Memory_45; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_175 = 6'h2e == L0Index ? io_FromL1 : L0Memory_46; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_176 = 6'h2f == L0Index ? io_FromL1 : L0Memory_47; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_177 = 6'h30 == L0Index ? io_FromL1 : L0Memory_48; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_178 = 6'h31 == L0Index ? io_FromL1 : L0Memory_49; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_179 = 6'h32 == L0Index ? io_FromL1 : L0Memory_50; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_180 = 6'h33 == L0Index ? io_FromL1 : L0Memory_51; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_181 = 6'h34 == L0Index ? io_FromL1 : L0Memory_52; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_182 = 6'h35 == L0Index ? io_FromL1 : L0Memory_53; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_183 = 6'h36 == L0Index ? io_FromL1 : L0Memory_54; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_184 = 6'h37 == L0Index ? io_FromL1 : L0Memory_55; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_185 = 6'h38 == L0Index ? io_FromL1 : L0Memory_56; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_186 = 6'h39 == L0Index ? io_FromL1 : L0Memory_57; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_187 = 6'h3a == L0Index ? io_FromL1 : L0Memory_58; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_188 = 6'h3b == L0Index ? io_FromL1 : L0Memory_59; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_189 = 6'h3c == L0Index ? io_FromL1 : L0Memory_60; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_190 = 6'h3d == L0Index ? io_FromL1 : L0Memory_61; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_191 = 6'h3e == L0Index ? io_FromL1 : L0Memory_62; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_192 = 6'h3f == L0Index ? io_FromL1 : L0Memory_63; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_193 = 7'h40 == _GEN_793 ? io_FromL1 : L0Memory_64; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_194 = 7'h41 == _GEN_793 ? io_FromL1 : L0Memory_65; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_195 = 7'h42 == _GEN_793 ? io_FromL1 : L0Memory_66; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_196 = 7'h43 == _GEN_793 ? io_FromL1 : L0Memory_67; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_197 = 7'h44 == _GEN_793 ? io_FromL1 : L0Memory_68; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_198 = 7'h45 == _GEN_793 ? io_FromL1 : L0Memory_69; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_199 = 7'h46 == _GEN_793 ? io_FromL1 : L0Memory_70; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_200 = 7'h47 == _GEN_793 ? io_FromL1 : L0Memory_71; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_201 = 7'h48 == _GEN_793 ? io_FromL1 : L0Memory_72; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_202 = 7'h49 == _GEN_793 ? io_FromL1 : L0Memory_73; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_203 = 7'h4a == _GEN_793 ? io_FromL1 : L0Memory_74; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_204 = 7'h4b == _GEN_793 ? io_FromL1 : L0Memory_75; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_205 = 7'h4c == _GEN_793 ? io_FromL1 : L0Memory_76; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_206 = 7'h4d == _GEN_793 ? io_FromL1 : L0Memory_77; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_207 = 7'h4e == _GEN_793 ? io_FromL1 : L0Memory_78; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_208 = 7'h4f == _GEN_793 ? io_FromL1 : L0Memory_79; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_209 = 7'h50 == _GEN_793 ? io_FromL1 : L0Memory_80; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_210 = 7'h51 == _GEN_793 ? io_FromL1 : L0Memory_81; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_211 = 7'h52 == _GEN_793 ? io_FromL1 : L0Memory_82; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_212 = 7'h53 == _GEN_793 ? io_FromL1 : L0Memory_83; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_213 = 7'h54 == _GEN_793 ? io_FromL1 : L0Memory_84; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_214 = 7'h55 == _GEN_793 ? io_FromL1 : L0Memory_85; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_215 = 7'h56 == _GEN_793 ? io_FromL1 : L0Memory_86; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_216 = 7'h57 == _GEN_793 ? io_FromL1 : L0Memory_87; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_217 = 7'h58 == _GEN_793 ? io_FromL1 : L0Memory_88; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_218 = 7'h59 == _GEN_793 ? io_FromL1 : L0Memory_89; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_219 = 7'h5a == _GEN_793 ? io_FromL1 : L0Memory_90; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_220 = 7'h5b == _GEN_793 ? io_FromL1 : L0Memory_91; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_221 = 7'h5c == _GEN_793 ? io_FromL1 : L0Memory_92; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_222 = 7'h5d == _GEN_793 ? io_FromL1 : L0Memory_93; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_223 = 7'h5e == _GEN_793 ? io_FromL1 : L0Memory_94; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_224 = 7'h5f == _GEN_793 ? io_FromL1 : L0Memory_95; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_225 = 7'h60 == _GEN_793 ? io_FromL1 : L0Memory_96; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_226 = 7'h61 == _GEN_793 ? io_FromL1 : L0Memory_97; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_227 = 7'h62 == _GEN_793 ? io_FromL1 : L0Memory_98; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_228 = 7'h63 == _GEN_793 ? io_FromL1 : L0Memory_99; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [5:0] _L0Index_T_2 = L0Index + 6'h1; // @[PEArray.scala 200:28]
  wire [15:0] _GEN_229 = count >= 10'h1 & count <= _T_27 ? _GEN_129 : L0Memory_0; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_230 = count >= 10'h1 & count <= _T_27 ? _GEN_130 : L0Memory_1; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_231 = count >= 10'h1 & count <= _T_27 ? _GEN_131 : L0Memory_2; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_232 = count >= 10'h1 & count <= _T_27 ? _GEN_132 : L0Memory_3; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_233 = count >= 10'h1 & count <= _T_27 ? _GEN_133 : L0Memory_4; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_234 = count >= 10'h1 & count <= _T_27 ? _GEN_134 : L0Memory_5; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_235 = count >= 10'h1 & count <= _T_27 ? _GEN_135 : L0Memory_6; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_236 = count >= 10'h1 & count <= _T_27 ? _GEN_136 : L0Memory_7; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_237 = count >= 10'h1 & count <= _T_27 ? _GEN_137 : L0Memory_8; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_238 = count >= 10'h1 & count <= _T_27 ? _GEN_138 : L0Memory_9; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_239 = count >= 10'h1 & count <= _T_27 ? _GEN_139 : L0Memory_10; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_240 = count >= 10'h1 & count <= _T_27 ? _GEN_140 : L0Memory_11; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_241 = count >= 10'h1 & count <= _T_27 ? _GEN_141 : L0Memory_12; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_242 = count >= 10'h1 & count <= _T_27 ? _GEN_142 : L0Memory_13; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_243 = count >= 10'h1 & count <= _T_27 ? _GEN_143 : L0Memory_14; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_244 = count >= 10'h1 & count <= _T_27 ? _GEN_144 : L0Memory_15; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_245 = count >= 10'h1 & count <= _T_27 ? _GEN_145 : L0Memory_16; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_246 = count >= 10'h1 & count <= _T_27 ? _GEN_146 : L0Memory_17; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_247 = count >= 10'h1 & count <= _T_27 ? _GEN_147 : L0Memory_18; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_248 = count >= 10'h1 & count <= _T_27 ? _GEN_148 : L0Memory_19; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_249 = count >= 10'h1 & count <= _T_27 ? _GEN_149 : L0Memory_20; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_250 = count >= 10'h1 & count <= _T_27 ? _GEN_150 : L0Memory_21; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_251 = count >= 10'h1 & count <= _T_27 ? _GEN_151 : L0Memory_22; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_252 = count >= 10'h1 & count <= _T_27 ? _GEN_152 : L0Memory_23; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_253 = count >= 10'h1 & count <= _T_27 ? _GEN_153 : L0Memory_24; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_254 = count >= 10'h1 & count <= _T_27 ? _GEN_154 : L0Memory_25; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_255 = count >= 10'h1 & count <= _T_27 ? _GEN_155 : L0Memory_26; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_256 = count >= 10'h1 & count <= _T_27 ? _GEN_156 : L0Memory_27; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_257 = count >= 10'h1 & count <= _T_27 ? _GEN_157 : L0Memory_28; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_258 = count >= 10'h1 & count <= _T_27 ? _GEN_158 : L0Memory_29; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_259 = count >= 10'h1 & count <= _T_27 ? _GEN_159 : L0Memory_30; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_260 = count >= 10'h1 & count <= _T_27 ? _GEN_160 : L0Memory_31; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_261 = count >= 10'h1 & count <= _T_27 ? _GEN_161 : L0Memory_32; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_262 = count >= 10'h1 & count <= _T_27 ? _GEN_162 : L0Memory_33; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_263 = count >= 10'h1 & count <= _T_27 ? _GEN_163 : L0Memory_34; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_264 = count >= 10'h1 & count <= _T_27 ? _GEN_164 : L0Memory_35; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_265 = count >= 10'h1 & count <= _T_27 ? _GEN_165 : L0Memory_36; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_266 = count >= 10'h1 & count <= _T_27 ? _GEN_166 : L0Memory_37; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_267 = count >= 10'h1 & count <= _T_27 ? _GEN_167 : L0Memory_38; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_268 = count >= 10'h1 & count <= _T_27 ? _GEN_168 : L0Memory_39; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_269 = count >= 10'h1 & count <= _T_27 ? _GEN_169 : L0Memory_40; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_270 = count >= 10'h1 & count <= _T_27 ? _GEN_170 : L0Memory_41; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_271 = count >= 10'h1 & count <= _T_27 ? _GEN_171 : L0Memory_42; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_272 = count >= 10'h1 & count <= _T_27 ? _GEN_172 : L0Memory_43; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_273 = count >= 10'h1 & count <= _T_27 ? _GEN_173 : L0Memory_44; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_274 = count >= 10'h1 & count <= _T_27 ? _GEN_174 : L0Memory_45; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_275 = count >= 10'h1 & count <= _T_27 ? _GEN_175 : L0Memory_46; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_276 = count >= 10'h1 & count <= _T_27 ? _GEN_176 : L0Memory_47; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_277 = count >= 10'h1 & count <= _T_27 ? _GEN_177 : L0Memory_48; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_278 = count >= 10'h1 & count <= _T_27 ? _GEN_178 : L0Memory_49; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_279 = count >= 10'h1 & count <= _T_27 ? _GEN_179 : L0Memory_50; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_280 = count >= 10'h1 & count <= _T_27 ? _GEN_180 : L0Memory_51; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_281 = count >= 10'h1 & count <= _T_27 ? _GEN_181 : L0Memory_52; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_282 = count >= 10'h1 & count <= _T_27 ? _GEN_182 : L0Memory_53; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_283 = count >= 10'h1 & count <= _T_27 ? _GEN_183 : L0Memory_54; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_284 = count >= 10'h1 & count <= _T_27 ? _GEN_184 : L0Memory_55; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_285 = count >= 10'h1 & count <= _T_27 ? _GEN_185 : L0Memory_56; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_286 = count >= 10'h1 & count <= _T_27 ? _GEN_186 : L0Memory_57; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_287 = count >= 10'h1 & count <= _T_27 ? _GEN_187 : L0Memory_58; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_288 = count >= 10'h1 & count <= _T_27 ? _GEN_188 : L0Memory_59; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_289 = count >= 10'h1 & count <= _T_27 ? _GEN_189 : L0Memory_60; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_290 = count >= 10'h1 & count <= _T_27 ? _GEN_190 : L0Memory_61; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_291 = count >= 10'h1 & count <= _T_27 ? _GEN_191 : L0Memory_62; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_292 = count >= 10'h1 & count <= _T_27 ? _GEN_192 : L0Memory_63; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_293 = count >= 10'h1 & count <= _T_27 ? _GEN_193 : L0Memory_64; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_294 = count >= 10'h1 & count <= _T_27 ? _GEN_194 : L0Memory_65; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_295 = count >= 10'h1 & count <= _T_27 ? _GEN_195 : L0Memory_66; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_296 = count >= 10'h1 & count <= _T_27 ? _GEN_196 : L0Memory_67; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_297 = count >= 10'h1 & count <= _T_27 ? _GEN_197 : L0Memory_68; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_298 = count >= 10'h1 & count <= _T_27 ? _GEN_198 : L0Memory_69; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_299 = count >= 10'h1 & count <= _T_27 ? _GEN_199 : L0Memory_70; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_300 = count >= 10'h1 & count <= _T_27 ? _GEN_200 : L0Memory_71; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_301 = count >= 10'h1 & count <= _T_27 ? _GEN_201 : L0Memory_72; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_302 = count >= 10'h1 & count <= _T_27 ? _GEN_202 : L0Memory_73; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_303 = count >= 10'h1 & count <= _T_27 ? _GEN_203 : L0Memory_74; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_304 = count >= 10'h1 & count <= _T_27 ? _GEN_204 : L0Memory_75; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_305 = count >= 10'h1 & count <= _T_27 ? _GEN_205 : L0Memory_76; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_306 = count >= 10'h1 & count <= _T_27 ? _GEN_206 : L0Memory_77; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_307 = count >= 10'h1 & count <= _T_27 ? _GEN_207 : L0Memory_78; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_308 = count >= 10'h1 & count <= _T_27 ? _GEN_208 : L0Memory_79; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_309 = count >= 10'h1 & count <= _T_27 ? _GEN_209 : L0Memory_80; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_310 = count >= 10'h1 & count <= _T_27 ? _GEN_210 : L0Memory_81; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_311 = count >= 10'h1 & count <= _T_27 ? _GEN_211 : L0Memory_82; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_312 = count >= 10'h1 & count <= _T_27 ? _GEN_212 : L0Memory_83; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_313 = count >= 10'h1 & count <= _T_27 ? _GEN_213 : L0Memory_84; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_314 = count >= 10'h1 & count <= _T_27 ? _GEN_214 : L0Memory_85; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_315 = count >= 10'h1 & count <= _T_27 ? _GEN_215 : L0Memory_86; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_316 = count >= 10'h1 & count <= _T_27 ? _GEN_216 : L0Memory_87; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_317 = count >= 10'h1 & count <= _T_27 ? _GEN_217 : L0Memory_88; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_318 = count >= 10'h1 & count <= _T_27 ? _GEN_218 : L0Memory_89; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_319 = count >= 10'h1 & count <= _T_27 ? _GEN_219 : L0Memory_90; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_320 = count >= 10'h1 & count <= _T_27 ? _GEN_220 : L0Memory_91; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_321 = count >= 10'h1 & count <= _T_27 ? _GEN_221 : L0Memory_92; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_322 = count >= 10'h1 & count <= _T_27 ? _GEN_222 : L0Memory_93; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_323 = count >= 10'h1 & count <= _T_27 ? _GEN_223 : L0Memory_94; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_324 = count >= 10'h1 & count <= _T_27 ? _GEN_224 : L0Memory_95; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_325 = count >= 10'h1 & count <= _T_27 ? _GEN_225 : L0Memory_96; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_326 = count >= 10'h1 & count <= _T_27 ? _GEN_226 : L0Memory_97; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_327 = count >= 10'h1 & count <= _T_27 ? _GEN_227 : L0Memory_98; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_328 = count >= 10'h1 & count <= _T_27 ? _GEN_228 : L0Memory_99; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [5:0] _GEN_329 = count >= 10'h1 & count <= _T_27 ? _L0Index_T_2 : _GEN_128; // @[PEArray.scala 198:59 PEArray.scala 200:17]
  wire [9:0] _GEN_330 = _T_24 ? 10'h0 : _GEN_127; // @[PEArray.scala 202:32 PEArray.scala 203:15]
  wire [2:0] _GEN_331 = _T_24 ? 3'h0 : state; // @[PEArray.scala 202:32 PEArray.scala 204:15 PEArray.scala 100:22]
  wire [9:0] _GEN_865 = {{4'd0}, GRU_out_width}; // @[PEArray.scala 220:19]
  wire [9:0] _GEN_0 = count % _GEN_865; // @[PEArray.scala 220:19]
  wire [5:0] _T_36 = _GEN_0[5:0]; // @[PEArray.scala 220:19]
  wire [5:0] _T_38 = GRU_out_width - 6'h1; // @[PEArray.scala 220:55]
  wire [5:0] _GEN_334 = _T_36 == _T_38 ? _L0Index_T_2 : 6'h0; // @[PEArray.scala 220:62 PEArray.scala 221:17 PEArray.scala 214:15]
  wire [5:0] _GEN_346 = _T_41 ? _GEN_334 : L0Index; // @[Conditional.scala 39:67 PEArray.scala 39:24]
  wire [9:0] _GEN_347 = _T_41 ? _GEN_330 : count; // @[Conditional.scala 39:67 PEArray.scala 101:22]
  wire [2:0] _GEN_348 = _T_41 ? _GEN_331 : state; // @[Conditional.scala 39:67 PEArray.scala 100:22]
  wire [5:0] _GEN_353 = _T_31 ? _GEN_334 : _GEN_346; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_354 = _T_31 ? _GEN_330 : _GEN_347; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_355 = _T_31 ? _GEN_331 : _GEN_348; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_356 = _T_22 ? _GEN_330 : _GEN_354; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_357 = _T_22 ? _GEN_329 : _GEN_353; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_458 = _T_22 ? _GEN_331 : _GEN_355; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_690 = _T_3 ? _GEN_118 : {{2'd0}, GRU_out_width}; // @[Conditional.scala 40:58 PEArray.scala 104:26]
  FP16MulAdder FP16MAC ( // @[PEArray.scala 72:23]
    .io_a(FP16MAC_io_a),
    .io_b(FP16MAC_io_b),
    .io_c(FP16MAC_io_c),
    .io_out(FP16MAC_io_out)
  );
  assign io_ToBelowPE = mux2out_reg; // @[PEArray.scala 94:16]
  assign FP16MAC_io_a = sel1 ? io_FromL1 : io_FromLeftPE; // @[PEArray.scala 50:14 PEArray.scala 50:23 PEArray.scala 51:24]
  assign FP16MAC_io_b = sel5 ? mux4out : _GEN_105; // @[PEArray.scala 77:13 PEArray.scala 78:18 PEArray.scala 81:18]
  assign FP16MAC_io_c = sel5 ? _GEN_105 : mux4out; // @[PEArray.scala 77:13 PEArray.scala 79:18 PEArray.scala 82:18]
  always @(posedge clock) begin
    if (reset) begin // @[PEArray.scala 39:24]
      L0Index <= 6'h0; // @[PEArray.scala 39:24]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h0; // @[PEArray.scala 159:15]
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        L0Index <= 6'he; // @[PEArray.scala 181:15]
      end else begin
        L0Index <= _GEN_357;
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_0 <= _GEN_229;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_1 <= _GEN_230;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_2 <= _GEN_231;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_3 <= _GEN_232;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_4 <= _GEN_233;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_5 <= _GEN_234;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_6 <= _GEN_235;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_7 <= _GEN_236;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_8 <= _GEN_237;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_9 <= _GEN_238;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_10 <= _GEN_239;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_11 <= _GEN_240;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_12 <= _GEN_241;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_13 <= _GEN_242;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_14 <= _GEN_243;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_15 <= _GEN_244;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_16 <= _GEN_245;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_17 <= _GEN_246;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_18 <= _GEN_247;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_19 <= _GEN_248;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_20 <= _GEN_249;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_21 <= _GEN_250;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_22 <= _GEN_251;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_23 <= _GEN_252;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_24 <= _GEN_253;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_25 <= _GEN_254;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_26 <= _GEN_255;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_27 <= _GEN_256;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_28 <= _GEN_257;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_29 <= _GEN_258;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_30 <= _GEN_259;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_31 <= _GEN_260;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_32 <= _GEN_261;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_33 <= _GEN_262;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_34 <= _GEN_263;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_35 <= _GEN_264;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_36 <= _GEN_265;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_37 <= _GEN_266;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_38 <= _GEN_267;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_39 <= _GEN_268;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_40 <= _GEN_269;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_41 <= _GEN_270;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_42 <= _GEN_271;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_43 <= _GEN_272;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_44 <= _GEN_273;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_45 <= _GEN_274;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_46 <= _GEN_275;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_47 <= _GEN_276;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_48 <= _GEN_277;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_49 <= _GEN_278;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_50 <= _GEN_279;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_51 <= _GEN_280;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_52 <= _GEN_281;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_53 <= _GEN_282;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_54 <= _GEN_283;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_55 <= _GEN_284;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_56 <= _GEN_285;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_57 <= _GEN_286;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_58 <= _GEN_287;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_59 <= _GEN_288;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_60 <= _GEN_289;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_61 <= _GEN_290;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_62 <= _GEN_291;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_63 <= _GEN_292;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_64 <= _GEN_293;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_65 <= _GEN_294;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_66 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_67 <= _GEN_296;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_68 <= _GEN_297;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_69 <= _GEN_298;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_70 <= _GEN_299;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_71 <= _GEN_300;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_72 <= _GEN_301;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_73 <= _GEN_302;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_74 <= _GEN_303;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_75 <= _GEN_304;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_76 <= _GEN_305;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_77 <= _GEN_306;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_78 <= _GEN_307;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_79 <= _GEN_308;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_80 <= _GEN_309;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_81 <= _GEN_310;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_82 <= _GEN_311;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_83 <= _GEN_312;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_84 <= _GEN_313;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_85 <= _GEN_314;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_86 <= _GEN_315;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_87 <= _GEN_316;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_88 <= _GEN_317;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_89 <= _GEN_318;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_90 <= _GEN_319;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_91 <= _GEN_320;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_92 <= _GEN_321;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_93 <= _GEN_322;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_94 <= _GEN_323;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_95 <= _GEN_324;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_96 <= _GEN_325;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_97 <= _GEN_326;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_98 <= _GEN_327;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_99 <= _GEN_328;
          end
        end
      end
    end
    if (reset) begin // @[PEArray.scala 100:22]
      state <= 3'h0; // @[PEArray.scala 100:22]
    end else if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[0]) begin // @[PEArray.scala 116:57]
        state <= 3'h1;
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      if (count == 10'h33) begin // @[PEArray.scala 164:27]
        state <= 3'h0; // @[PEArray.scala 166:15]
      end
    end else if (_T_16) begin // @[Conditional.scala 39:67]
      state <= _GEN_126;
    end else begin
      state <= _GEN_458;
    end
    if (reset) begin // @[PEArray.scala 90:28]
      mux2out_reg <= 16'h0; // @[PEArray.scala 90:28]
    end else begin
      mux2out_reg <= MAC_out; // @[PEArray.scala 90:28]
    end
    if (reset) begin // @[PEArray.scala 101:22]
      count <= 10'h0; // @[PEArray.scala 101:22]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        if (count == 10'h33) begin // @[PEArray.scala 164:27]
          count <= 10'h0; // @[PEArray.scala 165:15]
        end else begin
          count <= _GEN_120;
        end
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        count <= _GEN_125;
      end else begin
        count <= _GEN_356;
      end
    end
    GRU_out_width <= _GEN_690[5:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  L0Index = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  L0Memory_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  L0Memory_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  L0Memory_2 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  L0Memory_3 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  L0Memory_4 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  L0Memory_5 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  L0Memory_6 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  L0Memory_7 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  L0Memory_8 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  L0Memory_9 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  L0Memory_10 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  L0Memory_11 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  L0Memory_12 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  L0Memory_13 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  L0Memory_14 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  L0Memory_15 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  L0Memory_16 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  L0Memory_17 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  L0Memory_18 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  L0Memory_19 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  L0Memory_20 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  L0Memory_21 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  L0Memory_22 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  L0Memory_23 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  L0Memory_24 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  L0Memory_25 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  L0Memory_26 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  L0Memory_27 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  L0Memory_28 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  L0Memory_29 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  L0Memory_30 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  L0Memory_31 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  L0Memory_32 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  L0Memory_33 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  L0Memory_34 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  L0Memory_35 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  L0Memory_36 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  L0Memory_37 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  L0Memory_38 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  L0Memory_39 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  L0Memory_40 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  L0Memory_41 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  L0Memory_42 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  L0Memory_43 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  L0Memory_44 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  L0Memory_45 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  L0Memory_46 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  L0Memory_47 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  L0Memory_48 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  L0Memory_49 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  L0Memory_50 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  L0Memory_51 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  L0Memory_52 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  L0Memory_53 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  L0Memory_54 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  L0Memory_55 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  L0Memory_56 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  L0Memory_57 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  L0Memory_58 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  L0Memory_59 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  L0Memory_60 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  L0Memory_61 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  L0Memory_62 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  L0Memory_63 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  L0Memory_64 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  L0Memory_65 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  L0Memory_66 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  L0Memory_67 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  L0Memory_68 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  L0Memory_69 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  L0Memory_70 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  L0Memory_71 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  L0Memory_72 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  L0Memory_73 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  L0Memory_74 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  L0Memory_75 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  L0Memory_76 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  L0Memory_77 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  L0Memory_78 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  L0Memory_79 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  L0Memory_80 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  L0Memory_81 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  L0Memory_82 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  L0Memory_83 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  L0Memory_84 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  L0Memory_85 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  L0Memory_86 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  L0Memory_87 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  L0Memory_88 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  L0Memory_89 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  L0Memory_90 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  L0Memory_91 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  L0Memory_92 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  L0Memory_93 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  L0Memory_94 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  L0Memory_95 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  L0Memory_96 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  L0Memory_97 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  L0Memory_98 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  L0Memory_99 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  state = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  mux2out_reg = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  count = _RAND_103[9:0];
  _RAND_104 = {1{`RANDOM}};
  GRU_out_width = _RAND_104[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PE_34(
  input         clock,
  input         reset,
  input  [15:0] io_FromAbovePE,
  input  [15:0] io_FromLeftPE,
  input  [15:0] io_FromL1,
  input  [11:0] io_control_signal_mask,
  output [15:0] io_ToBelowPE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] FP16MAC_io_a; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_b; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_c; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_out; // @[PEArray.scala 72:23]
  reg [5:0] L0Index; // @[PEArray.scala 39:24]
  reg [15:0] L0Memory_0; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_1; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_2; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_3; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_4; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_5; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_6; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_7; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_8; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_9; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_10; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_11; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_12; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_13; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_14; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_15; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_16; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_17; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_18; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_19; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_20; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_21; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_22; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_23; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_24; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_25; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_26; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_27; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_28; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_29; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_30; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_31; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_32; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_33; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_34; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_35; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_36; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_37; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_38; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_39; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_40; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_41; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_42; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_43; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_44; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_45; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_46; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_47; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_48; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_49; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_50; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_51; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_52; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_53; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_54; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_55; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_56; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_57; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_58; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_59; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_60; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_61; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_62; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_63; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_64; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_65; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_66; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_67; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_68; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_69; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_70; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_71; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_72; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_73; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_74; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_75; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_76; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_77; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_78; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_79; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_80; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_81; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_82; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_83; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_84; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_85; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_86; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_87; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_88; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_89; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_90; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_91; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_92; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_93; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_94; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_95; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_96; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_97; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_98; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_99; // @[PEArray.scala 40:21]
  reg [2:0] state; // @[PEArray.scala 100:22]
  wire  _T_3 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_12 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_16 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_22 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_31 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_41 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_342 = _T_41 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 231:12 PEArray.scala 32:8]
  wire  _GEN_349 = _T_31 ? 1'h0 : _GEN_342; // @[Conditional.scala 39:67 PEArray.scala 208:12]
  wire  _GEN_459 = _T_22 | _GEN_349; // @[Conditional.scala 39:67 PEArray.scala 32:8]
  wire  _GEN_463 = _T_16 ? 1'h0 : _GEN_459; // @[Conditional.scala 39:67]
  wire  _GEN_572 = _T_12 | _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 149:12]
  wire  sel1 = _T_3 | _GEN_572; // @[Conditional.scala 40:58 PEArray.scala 108:12]
  wire [15:0] MAC_out = FP16MAC_io_out; // @[PEArray.scala 47:21 PEArray.scala 85:11]
  wire [1:0] _GEN_344 = _T_41 ? 2'h2 : 2'h0; // @[Conditional.scala 39:67 PEArray.scala 233:12 PEArray.scala 35:8]
  wire [1:0] _GEN_351 = _T_31 ? 2'h2 : _GEN_344; // @[Conditional.scala 39:67 PEArray.scala 210:12]
  wire [1:0] _GEN_461 = _T_22 ? 2'h0 : _GEN_351; // @[Conditional.scala 39:67 PEArray.scala 35:8]
  wire [1:0] _GEN_466 = _T_16 ? 2'h0 : _GEN_461; // @[Conditional.scala 39:67 PEArray.scala 178:12]
  wire [1:0] _GEN_574 = _T_12 ? 2'h1 : _GEN_466; // @[Conditional.scala 39:67]
  wire [1:0] sel4 = _T_3 ? 2'h0 : _GEN_574; // @[Conditional.scala 40:58 PEArray.scala 111:12]
  wire [15:0] _GEN_3 = sel4 == 2'h2 ? io_FromL1 : 16'h0; // @[PEArray.scala 65:28 PEArray.scala 66:15 PEArray.scala 69:15]
  wire [15:0] _GEN_4 = sel4 == 2'h1 ? io_FromAbovePE : _GEN_3; // @[PEArray.scala 62:28 PEArray.scala 63:15]
  wire [15:0] mux4out = sel4 == 2'h0 ? 16'h0 : _GEN_4; // @[PEArray.scala 59:22 PEArray.scala 60:13]
  wire [15:0] _GEN_7 = 6'h1 == L0Index ? L0Memory_1 : L0Memory_0; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_8 = 6'h2 == L0Index ? L0Memory_2 : _GEN_7; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_9 = 6'h3 == L0Index ? L0Memory_3 : _GEN_8; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_10 = 6'h4 == L0Index ? L0Memory_4 : _GEN_9; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_11 = 6'h5 == L0Index ? L0Memory_5 : _GEN_10; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_12 = 6'h6 == L0Index ? L0Memory_6 : _GEN_11; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_13 = 6'h7 == L0Index ? L0Memory_7 : _GEN_12; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_14 = 6'h8 == L0Index ? L0Memory_8 : _GEN_13; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_15 = 6'h9 == L0Index ? L0Memory_9 : _GEN_14; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_16 = 6'ha == L0Index ? L0Memory_10 : _GEN_15; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_17 = 6'hb == L0Index ? L0Memory_11 : _GEN_16; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_18 = 6'hc == L0Index ? L0Memory_12 : _GEN_17; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_19 = 6'hd == L0Index ? L0Memory_13 : _GEN_18; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_20 = 6'he == L0Index ? L0Memory_14 : _GEN_19; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_21 = 6'hf == L0Index ? L0Memory_15 : _GEN_20; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_22 = 6'h10 == L0Index ? L0Memory_16 : _GEN_21; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_23 = 6'h11 == L0Index ? L0Memory_17 : _GEN_22; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_24 = 6'h12 == L0Index ? L0Memory_18 : _GEN_23; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_25 = 6'h13 == L0Index ? L0Memory_19 : _GEN_24; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_26 = 6'h14 == L0Index ? L0Memory_20 : _GEN_25; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_27 = 6'h15 == L0Index ? L0Memory_21 : _GEN_26; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_28 = 6'h16 == L0Index ? L0Memory_22 : _GEN_27; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_29 = 6'h17 == L0Index ? L0Memory_23 : _GEN_28; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_30 = 6'h18 == L0Index ? L0Memory_24 : _GEN_29; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_31 = 6'h19 == L0Index ? L0Memory_25 : _GEN_30; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_32 = 6'h1a == L0Index ? L0Memory_26 : _GEN_31; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_33 = 6'h1b == L0Index ? L0Memory_27 : _GEN_32; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_34 = 6'h1c == L0Index ? L0Memory_28 : _GEN_33; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_35 = 6'h1d == L0Index ? L0Memory_29 : _GEN_34; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_36 = 6'h1e == L0Index ? L0Memory_30 : _GEN_35; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_37 = 6'h1f == L0Index ? L0Memory_31 : _GEN_36; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_38 = 6'h20 == L0Index ? L0Memory_32 : _GEN_37; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_39 = 6'h21 == L0Index ? L0Memory_33 : _GEN_38; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_40 = 6'h22 == L0Index ? L0Memory_34 : _GEN_39; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_41 = 6'h23 == L0Index ? L0Memory_35 : _GEN_40; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_42 = 6'h24 == L0Index ? L0Memory_36 : _GEN_41; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_43 = 6'h25 == L0Index ? L0Memory_37 : _GEN_42; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_44 = 6'h26 == L0Index ? L0Memory_38 : _GEN_43; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_45 = 6'h27 == L0Index ? L0Memory_39 : _GEN_44; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_46 = 6'h28 == L0Index ? L0Memory_40 : _GEN_45; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_47 = 6'h29 == L0Index ? L0Memory_41 : _GEN_46; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_48 = 6'h2a == L0Index ? L0Memory_42 : _GEN_47; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_49 = 6'h2b == L0Index ? L0Memory_43 : _GEN_48; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_50 = 6'h2c == L0Index ? L0Memory_44 : _GEN_49; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_51 = 6'h2d == L0Index ? L0Memory_45 : _GEN_50; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_52 = 6'h2e == L0Index ? L0Memory_46 : _GEN_51; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_53 = 6'h2f == L0Index ? L0Memory_47 : _GEN_52; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_54 = 6'h30 == L0Index ? L0Memory_48 : _GEN_53; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_55 = 6'h31 == L0Index ? L0Memory_49 : _GEN_54; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_56 = 6'h32 == L0Index ? L0Memory_50 : _GEN_55; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_57 = 6'h33 == L0Index ? L0Memory_51 : _GEN_56; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_58 = 6'h34 == L0Index ? L0Memory_52 : _GEN_57; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_59 = 6'h35 == L0Index ? L0Memory_53 : _GEN_58; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_60 = 6'h36 == L0Index ? L0Memory_54 : _GEN_59; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_61 = 6'h37 == L0Index ? L0Memory_55 : _GEN_60; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_62 = 6'h38 == L0Index ? L0Memory_56 : _GEN_61; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_63 = 6'h39 == L0Index ? L0Memory_57 : _GEN_62; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_64 = 6'h3a == L0Index ? L0Memory_58 : _GEN_63; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_65 = 6'h3b == L0Index ? L0Memory_59 : _GEN_64; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_66 = 6'h3c == L0Index ? L0Memory_60 : _GEN_65; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_67 = 6'h3d == L0Index ? L0Memory_61 : _GEN_66; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_68 = 6'h3e == L0Index ? L0Memory_62 : _GEN_67; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_69 = 6'h3f == L0Index ? L0Memory_63 : _GEN_68; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [6:0] _GEN_793 = {{1'd0}, L0Index}; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_70 = 7'h40 == _GEN_793 ? L0Memory_64 : _GEN_69; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_71 = 7'h41 == _GEN_793 ? L0Memory_65 : _GEN_70; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_72 = 7'h42 == _GEN_793 ? L0Memory_66 : _GEN_71; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_73 = 7'h43 == _GEN_793 ? L0Memory_67 : _GEN_72; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_74 = 7'h44 == _GEN_793 ? L0Memory_68 : _GEN_73; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_75 = 7'h45 == _GEN_793 ? L0Memory_69 : _GEN_74; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_76 = 7'h46 == _GEN_793 ? L0Memory_70 : _GEN_75; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_77 = 7'h47 == _GEN_793 ? L0Memory_71 : _GEN_76; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_78 = 7'h48 == _GEN_793 ? L0Memory_72 : _GEN_77; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_79 = 7'h49 == _GEN_793 ? L0Memory_73 : _GEN_78; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_80 = 7'h4a == _GEN_793 ? L0Memory_74 : _GEN_79; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_81 = 7'h4b == _GEN_793 ? L0Memory_75 : _GEN_80; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_82 = 7'h4c == _GEN_793 ? L0Memory_76 : _GEN_81; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_83 = 7'h4d == _GEN_793 ? L0Memory_77 : _GEN_82; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_84 = 7'h4e == _GEN_793 ? L0Memory_78 : _GEN_83; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_85 = 7'h4f == _GEN_793 ? L0Memory_79 : _GEN_84; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_86 = 7'h50 == _GEN_793 ? L0Memory_80 : _GEN_85; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_87 = 7'h51 == _GEN_793 ? L0Memory_81 : _GEN_86; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_88 = 7'h52 == _GEN_793 ? L0Memory_82 : _GEN_87; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_89 = 7'h53 == _GEN_793 ? L0Memory_83 : _GEN_88; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_90 = 7'h54 == _GEN_793 ? L0Memory_84 : _GEN_89; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_91 = 7'h55 == _GEN_793 ? L0Memory_85 : _GEN_90; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_92 = 7'h56 == _GEN_793 ? L0Memory_86 : _GEN_91; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_93 = 7'h57 == _GEN_793 ? L0Memory_87 : _GEN_92; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_94 = 7'h58 == _GEN_793 ? L0Memory_88 : _GEN_93; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_95 = 7'h59 == _GEN_793 ? L0Memory_89 : _GEN_94; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_96 = 7'h5a == _GEN_793 ? L0Memory_90 : _GEN_95; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_97 = 7'h5b == _GEN_793 ? L0Memory_91 : _GEN_96; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_98 = 7'h5c == _GEN_793 ? L0Memory_92 : _GEN_97; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_99 = 7'h5d == _GEN_793 ? L0Memory_93 : _GEN_98; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_100 = 7'h5e == _GEN_793 ? L0Memory_94 : _GEN_99; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_101 = 7'h5f == _GEN_793 ? L0Memory_95 : _GEN_100; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_102 = 7'h60 == _GEN_793 ? L0Memory_96 : _GEN_101; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_103 = 7'h61 == _GEN_793 ? L0Memory_97 : _GEN_102; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_104 = 7'h62 == _GEN_793 ? L0Memory_98 : _GEN_103; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_105 = 7'h63 == _GEN_793 ? L0Memory_99 : _GEN_104; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire  _GEN_575 = _T_12 ? 1'h0 : _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 157:12]
  wire  sel5 = _T_3 ? 1'h0 : _GEN_575; // @[Conditional.scala 40:58 PEArray.scala 112:12]
  reg [15:0] mux2out_reg; // @[PEArray.scala 90:28]
  reg [9:0] count; // @[PEArray.scala 101:22]
  reg [5:0] GRU_out_width; // @[PEArray.scala 104:26]
  wire [7:0] _GEN_118 = io_control_signal_mask[0] ? 8'h0 : {{2'd0}, GRU_out_width}; // @[PEArray.scala 116:57 PEArray.scala 145:23 PEArray.scala 104:26]
  wire [9:0] _count_T_1 = count + 10'h1; // @[PEArray.scala 162:24]
  wire [9:0] _GEN_120 = count != 10'h33 ? _count_T_1 : count; // @[PEArray.scala 161:27 PEArray.scala 162:15 PEArray.scala 101:22]
  wire [9:0] _GEN_124 = count != 10'h188 ? _count_T_1 : count; // @[PEArray.scala 183:28 PEArray.scala 184:15 PEArray.scala 101:22]
  wire [9:0] _GEN_125 = count == 10'h188 ? 10'h0 : _GEN_124; // @[PEArray.scala 186:28 PEArray.scala 187:15]
  wire [2:0] _GEN_126 = count == 10'h188 ? 3'h0 : state; // @[PEArray.scala 186:28 PEArray.scala 188:15 PEArray.scala 100:22]
  wire [9:0] _GEN_127 = count != 10'h0 ? _count_T_1 : count; // @[PEArray.scala 192:32 PEArray.scala 193:15 PEArray.scala 101:22]
  wire  _T_24 = count == 10'h0; // @[PEArray.scala 195:18]
  wire [5:0] _GEN_128 = count == 10'h0 ? 6'h0 : L0Index; // @[PEArray.scala 195:26 PEArray.scala 196:17 PEArray.scala 39:24]
  wire [9:0] _T_27 = 10'h0 - 10'h1; // @[PEArray.scala 198:51]
  wire [15:0] _GEN_129 = 6'h0 == L0Index ? io_FromL1 : L0Memory_0; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_130 = 6'h1 == L0Index ? io_FromL1 : L0Memory_1; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_131 = 6'h2 == L0Index ? io_FromL1 : L0Memory_2; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_132 = 6'h3 == L0Index ? io_FromL1 : L0Memory_3; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_133 = 6'h4 == L0Index ? io_FromL1 : L0Memory_4; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_134 = 6'h5 == L0Index ? io_FromL1 : L0Memory_5; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_135 = 6'h6 == L0Index ? io_FromL1 : L0Memory_6; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_136 = 6'h7 == L0Index ? io_FromL1 : L0Memory_7; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_137 = 6'h8 == L0Index ? io_FromL1 : L0Memory_8; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_138 = 6'h9 == L0Index ? io_FromL1 : L0Memory_9; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_139 = 6'ha == L0Index ? io_FromL1 : L0Memory_10; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_140 = 6'hb == L0Index ? io_FromL1 : L0Memory_11; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_141 = 6'hc == L0Index ? io_FromL1 : L0Memory_12; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_142 = 6'hd == L0Index ? io_FromL1 : L0Memory_13; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_143 = 6'he == L0Index ? io_FromL1 : L0Memory_14; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_144 = 6'hf == L0Index ? io_FromL1 : L0Memory_15; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_145 = 6'h10 == L0Index ? io_FromL1 : L0Memory_16; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_146 = 6'h11 == L0Index ? io_FromL1 : L0Memory_17; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_147 = 6'h12 == L0Index ? io_FromL1 : L0Memory_18; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_148 = 6'h13 == L0Index ? io_FromL1 : L0Memory_19; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_149 = 6'h14 == L0Index ? io_FromL1 : L0Memory_20; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_150 = 6'h15 == L0Index ? io_FromL1 : L0Memory_21; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_151 = 6'h16 == L0Index ? io_FromL1 : L0Memory_22; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_152 = 6'h17 == L0Index ? io_FromL1 : L0Memory_23; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_153 = 6'h18 == L0Index ? io_FromL1 : L0Memory_24; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_154 = 6'h19 == L0Index ? io_FromL1 : L0Memory_25; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_155 = 6'h1a == L0Index ? io_FromL1 : L0Memory_26; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_156 = 6'h1b == L0Index ? io_FromL1 : L0Memory_27; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_157 = 6'h1c == L0Index ? io_FromL1 : L0Memory_28; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_158 = 6'h1d == L0Index ? io_FromL1 : L0Memory_29; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_159 = 6'h1e == L0Index ? io_FromL1 : L0Memory_30; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_160 = 6'h1f == L0Index ? io_FromL1 : L0Memory_31; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_161 = 6'h20 == L0Index ? io_FromL1 : L0Memory_32; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_162 = 6'h21 == L0Index ? io_FromL1 : L0Memory_33; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_163 = 6'h22 == L0Index ? io_FromL1 : L0Memory_34; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_164 = 6'h23 == L0Index ? io_FromL1 : L0Memory_35; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_165 = 6'h24 == L0Index ? io_FromL1 : L0Memory_36; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_166 = 6'h25 == L0Index ? io_FromL1 : L0Memory_37; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_167 = 6'h26 == L0Index ? io_FromL1 : L0Memory_38; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_168 = 6'h27 == L0Index ? io_FromL1 : L0Memory_39; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_169 = 6'h28 == L0Index ? io_FromL1 : L0Memory_40; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_170 = 6'h29 == L0Index ? io_FromL1 : L0Memory_41; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_171 = 6'h2a == L0Index ? io_FromL1 : L0Memory_42; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_172 = 6'h2b == L0Index ? io_FromL1 : L0Memory_43; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_173 = 6'h2c == L0Index ? io_FromL1 : L0Memory_44; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_174 = 6'h2d == L0Index ? io_FromL1 : L0Memory_45; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_175 = 6'h2e == L0Index ? io_FromL1 : L0Memory_46; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_176 = 6'h2f == L0Index ? io_FromL1 : L0Memory_47; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_177 = 6'h30 == L0Index ? io_FromL1 : L0Memory_48; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_178 = 6'h31 == L0Index ? io_FromL1 : L0Memory_49; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_179 = 6'h32 == L0Index ? io_FromL1 : L0Memory_50; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_180 = 6'h33 == L0Index ? io_FromL1 : L0Memory_51; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_181 = 6'h34 == L0Index ? io_FromL1 : L0Memory_52; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_182 = 6'h35 == L0Index ? io_FromL1 : L0Memory_53; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_183 = 6'h36 == L0Index ? io_FromL1 : L0Memory_54; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_184 = 6'h37 == L0Index ? io_FromL1 : L0Memory_55; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_185 = 6'h38 == L0Index ? io_FromL1 : L0Memory_56; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_186 = 6'h39 == L0Index ? io_FromL1 : L0Memory_57; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_187 = 6'h3a == L0Index ? io_FromL1 : L0Memory_58; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_188 = 6'h3b == L0Index ? io_FromL1 : L0Memory_59; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_189 = 6'h3c == L0Index ? io_FromL1 : L0Memory_60; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_190 = 6'h3d == L0Index ? io_FromL1 : L0Memory_61; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_191 = 6'h3e == L0Index ? io_FromL1 : L0Memory_62; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_192 = 6'h3f == L0Index ? io_FromL1 : L0Memory_63; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_193 = 7'h40 == _GEN_793 ? io_FromL1 : L0Memory_64; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_194 = 7'h41 == _GEN_793 ? io_FromL1 : L0Memory_65; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_195 = 7'h42 == _GEN_793 ? io_FromL1 : L0Memory_66; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_196 = 7'h43 == _GEN_793 ? io_FromL1 : L0Memory_67; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_197 = 7'h44 == _GEN_793 ? io_FromL1 : L0Memory_68; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_198 = 7'h45 == _GEN_793 ? io_FromL1 : L0Memory_69; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_199 = 7'h46 == _GEN_793 ? io_FromL1 : L0Memory_70; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_200 = 7'h47 == _GEN_793 ? io_FromL1 : L0Memory_71; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_201 = 7'h48 == _GEN_793 ? io_FromL1 : L0Memory_72; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_202 = 7'h49 == _GEN_793 ? io_FromL1 : L0Memory_73; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_203 = 7'h4a == _GEN_793 ? io_FromL1 : L0Memory_74; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_204 = 7'h4b == _GEN_793 ? io_FromL1 : L0Memory_75; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_205 = 7'h4c == _GEN_793 ? io_FromL1 : L0Memory_76; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_206 = 7'h4d == _GEN_793 ? io_FromL1 : L0Memory_77; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_207 = 7'h4e == _GEN_793 ? io_FromL1 : L0Memory_78; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_208 = 7'h4f == _GEN_793 ? io_FromL1 : L0Memory_79; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_209 = 7'h50 == _GEN_793 ? io_FromL1 : L0Memory_80; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_210 = 7'h51 == _GEN_793 ? io_FromL1 : L0Memory_81; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_211 = 7'h52 == _GEN_793 ? io_FromL1 : L0Memory_82; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_212 = 7'h53 == _GEN_793 ? io_FromL1 : L0Memory_83; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_213 = 7'h54 == _GEN_793 ? io_FromL1 : L0Memory_84; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_214 = 7'h55 == _GEN_793 ? io_FromL1 : L0Memory_85; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_215 = 7'h56 == _GEN_793 ? io_FromL1 : L0Memory_86; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_216 = 7'h57 == _GEN_793 ? io_FromL1 : L0Memory_87; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_217 = 7'h58 == _GEN_793 ? io_FromL1 : L0Memory_88; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_218 = 7'h59 == _GEN_793 ? io_FromL1 : L0Memory_89; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_219 = 7'h5a == _GEN_793 ? io_FromL1 : L0Memory_90; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_220 = 7'h5b == _GEN_793 ? io_FromL1 : L0Memory_91; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_221 = 7'h5c == _GEN_793 ? io_FromL1 : L0Memory_92; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_222 = 7'h5d == _GEN_793 ? io_FromL1 : L0Memory_93; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_223 = 7'h5e == _GEN_793 ? io_FromL1 : L0Memory_94; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_224 = 7'h5f == _GEN_793 ? io_FromL1 : L0Memory_95; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_225 = 7'h60 == _GEN_793 ? io_FromL1 : L0Memory_96; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_226 = 7'h61 == _GEN_793 ? io_FromL1 : L0Memory_97; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_227 = 7'h62 == _GEN_793 ? io_FromL1 : L0Memory_98; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_228 = 7'h63 == _GEN_793 ? io_FromL1 : L0Memory_99; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [5:0] _L0Index_T_2 = L0Index + 6'h1; // @[PEArray.scala 200:28]
  wire [15:0] _GEN_229 = count >= 10'h1 & count <= _T_27 ? _GEN_129 : L0Memory_0; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_230 = count >= 10'h1 & count <= _T_27 ? _GEN_130 : L0Memory_1; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_231 = count >= 10'h1 & count <= _T_27 ? _GEN_131 : L0Memory_2; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_232 = count >= 10'h1 & count <= _T_27 ? _GEN_132 : L0Memory_3; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_233 = count >= 10'h1 & count <= _T_27 ? _GEN_133 : L0Memory_4; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_234 = count >= 10'h1 & count <= _T_27 ? _GEN_134 : L0Memory_5; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_235 = count >= 10'h1 & count <= _T_27 ? _GEN_135 : L0Memory_6; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_236 = count >= 10'h1 & count <= _T_27 ? _GEN_136 : L0Memory_7; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_237 = count >= 10'h1 & count <= _T_27 ? _GEN_137 : L0Memory_8; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_238 = count >= 10'h1 & count <= _T_27 ? _GEN_138 : L0Memory_9; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_239 = count >= 10'h1 & count <= _T_27 ? _GEN_139 : L0Memory_10; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_240 = count >= 10'h1 & count <= _T_27 ? _GEN_140 : L0Memory_11; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_241 = count >= 10'h1 & count <= _T_27 ? _GEN_141 : L0Memory_12; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_242 = count >= 10'h1 & count <= _T_27 ? _GEN_142 : L0Memory_13; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_243 = count >= 10'h1 & count <= _T_27 ? _GEN_143 : L0Memory_14; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_244 = count >= 10'h1 & count <= _T_27 ? _GEN_144 : L0Memory_15; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_245 = count >= 10'h1 & count <= _T_27 ? _GEN_145 : L0Memory_16; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_246 = count >= 10'h1 & count <= _T_27 ? _GEN_146 : L0Memory_17; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_247 = count >= 10'h1 & count <= _T_27 ? _GEN_147 : L0Memory_18; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_248 = count >= 10'h1 & count <= _T_27 ? _GEN_148 : L0Memory_19; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_249 = count >= 10'h1 & count <= _T_27 ? _GEN_149 : L0Memory_20; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_250 = count >= 10'h1 & count <= _T_27 ? _GEN_150 : L0Memory_21; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_251 = count >= 10'h1 & count <= _T_27 ? _GEN_151 : L0Memory_22; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_252 = count >= 10'h1 & count <= _T_27 ? _GEN_152 : L0Memory_23; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_253 = count >= 10'h1 & count <= _T_27 ? _GEN_153 : L0Memory_24; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_254 = count >= 10'h1 & count <= _T_27 ? _GEN_154 : L0Memory_25; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_255 = count >= 10'h1 & count <= _T_27 ? _GEN_155 : L0Memory_26; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_256 = count >= 10'h1 & count <= _T_27 ? _GEN_156 : L0Memory_27; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_257 = count >= 10'h1 & count <= _T_27 ? _GEN_157 : L0Memory_28; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_258 = count >= 10'h1 & count <= _T_27 ? _GEN_158 : L0Memory_29; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_259 = count >= 10'h1 & count <= _T_27 ? _GEN_159 : L0Memory_30; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_260 = count >= 10'h1 & count <= _T_27 ? _GEN_160 : L0Memory_31; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_261 = count >= 10'h1 & count <= _T_27 ? _GEN_161 : L0Memory_32; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_262 = count >= 10'h1 & count <= _T_27 ? _GEN_162 : L0Memory_33; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_263 = count >= 10'h1 & count <= _T_27 ? _GEN_163 : L0Memory_34; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_264 = count >= 10'h1 & count <= _T_27 ? _GEN_164 : L0Memory_35; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_265 = count >= 10'h1 & count <= _T_27 ? _GEN_165 : L0Memory_36; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_266 = count >= 10'h1 & count <= _T_27 ? _GEN_166 : L0Memory_37; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_267 = count >= 10'h1 & count <= _T_27 ? _GEN_167 : L0Memory_38; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_268 = count >= 10'h1 & count <= _T_27 ? _GEN_168 : L0Memory_39; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_269 = count >= 10'h1 & count <= _T_27 ? _GEN_169 : L0Memory_40; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_270 = count >= 10'h1 & count <= _T_27 ? _GEN_170 : L0Memory_41; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_271 = count >= 10'h1 & count <= _T_27 ? _GEN_171 : L0Memory_42; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_272 = count >= 10'h1 & count <= _T_27 ? _GEN_172 : L0Memory_43; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_273 = count >= 10'h1 & count <= _T_27 ? _GEN_173 : L0Memory_44; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_274 = count >= 10'h1 & count <= _T_27 ? _GEN_174 : L0Memory_45; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_275 = count >= 10'h1 & count <= _T_27 ? _GEN_175 : L0Memory_46; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_276 = count >= 10'h1 & count <= _T_27 ? _GEN_176 : L0Memory_47; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_277 = count >= 10'h1 & count <= _T_27 ? _GEN_177 : L0Memory_48; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_278 = count >= 10'h1 & count <= _T_27 ? _GEN_178 : L0Memory_49; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_279 = count >= 10'h1 & count <= _T_27 ? _GEN_179 : L0Memory_50; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_280 = count >= 10'h1 & count <= _T_27 ? _GEN_180 : L0Memory_51; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_281 = count >= 10'h1 & count <= _T_27 ? _GEN_181 : L0Memory_52; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_282 = count >= 10'h1 & count <= _T_27 ? _GEN_182 : L0Memory_53; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_283 = count >= 10'h1 & count <= _T_27 ? _GEN_183 : L0Memory_54; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_284 = count >= 10'h1 & count <= _T_27 ? _GEN_184 : L0Memory_55; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_285 = count >= 10'h1 & count <= _T_27 ? _GEN_185 : L0Memory_56; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_286 = count >= 10'h1 & count <= _T_27 ? _GEN_186 : L0Memory_57; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_287 = count >= 10'h1 & count <= _T_27 ? _GEN_187 : L0Memory_58; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_288 = count >= 10'h1 & count <= _T_27 ? _GEN_188 : L0Memory_59; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_289 = count >= 10'h1 & count <= _T_27 ? _GEN_189 : L0Memory_60; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_290 = count >= 10'h1 & count <= _T_27 ? _GEN_190 : L0Memory_61; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_291 = count >= 10'h1 & count <= _T_27 ? _GEN_191 : L0Memory_62; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_292 = count >= 10'h1 & count <= _T_27 ? _GEN_192 : L0Memory_63; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_293 = count >= 10'h1 & count <= _T_27 ? _GEN_193 : L0Memory_64; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_294 = count >= 10'h1 & count <= _T_27 ? _GEN_194 : L0Memory_65; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_295 = count >= 10'h1 & count <= _T_27 ? _GEN_195 : L0Memory_66; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_296 = count >= 10'h1 & count <= _T_27 ? _GEN_196 : L0Memory_67; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_297 = count >= 10'h1 & count <= _T_27 ? _GEN_197 : L0Memory_68; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_298 = count >= 10'h1 & count <= _T_27 ? _GEN_198 : L0Memory_69; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_299 = count >= 10'h1 & count <= _T_27 ? _GEN_199 : L0Memory_70; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_300 = count >= 10'h1 & count <= _T_27 ? _GEN_200 : L0Memory_71; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_301 = count >= 10'h1 & count <= _T_27 ? _GEN_201 : L0Memory_72; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_302 = count >= 10'h1 & count <= _T_27 ? _GEN_202 : L0Memory_73; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_303 = count >= 10'h1 & count <= _T_27 ? _GEN_203 : L0Memory_74; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_304 = count >= 10'h1 & count <= _T_27 ? _GEN_204 : L0Memory_75; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_305 = count >= 10'h1 & count <= _T_27 ? _GEN_205 : L0Memory_76; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_306 = count >= 10'h1 & count <= _T_27 ? _GEN_206 : L0Memory_77; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_307 = count >= 10'h1 & count <= _T_27 ? _GEN_207 : L0Memory_78; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_308 = count >= 10'h1 & count <= _T_27 ? _GEN_208 : L0Memory_79; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_309 = count >= 10'h1 & count <= _T_27 ? _GEN_209 : L0Memory_80; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_310 = count >= 10'h1 & count <= _T_27 ? _GEN_210 : L0Memory_81; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_311 = count >= 10'h1 & count <= _T_27 ? _GEN_211 : L0Memory_82; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_312 = count >= 10'h1 & count <= _T_27 ? _GEN_212 : L0Memory_83; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_313 = count >= 10'h1 & count <= _T_27 ? _GEN_213 : L0Memory_84; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_314 = count >= 10'h1 & count <= _T_27 ? _GEN_214 : L0Memory_85; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_315 = count >= 10'h1 & count <= _T_27 ? _GEN_215 : L0Memory_86; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_316 = count >= 10'h1 & count <= _T_27 ? _GEN_216 : L0Memory_87; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_317 = count >= 10'h1 & count <= _T_27 ? _GEN_217 : L0Memory_88; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_318 = count >= 10'h1 & count <= _T_27 ? _GEN_218 : L0Memory_89; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_319 = count >= 10'h1 & count <= _T_27 ? _GEN_219 : L0Memory_90; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_320 = count >= 10'h1 & count <= _T_27 ? _GEN_220 : L0Memory_91; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_321 = count >= 10'h1 & count <= _T_27 ? _GEN_221 : L0Memory_92; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_322 = count >= 10'h1 & count <= _T_27 ? _GEN_222 : L0Memory_93; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_323 = count >= 10'h1 & count <= _T_27 ? _GEN_223 : L0Memory_94; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_324 = count >= 10'h1 & count <= _T_27 ? _GEN_224 : L0Memory_95; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_325 = count >= 10'h1 & count <= _T_27 ? _GEN_225 : L0Memory_96; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_326 = count >= 10'h1 & count <= _T_27 ? _GEN_226 : L0Memory_97; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_327 = count >= 10'h1 & count <= _T_27 ? _GEN_227 : L0Memory_98; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_328 = count >= 10'h1 & count <= _T_27 ? _GEN_228 : L0Memory_99; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [5:0] _GEN_329 = count >= 10'h1 & count <= _T_27 ? _L0Index_T_2 : _GEN_128; // @[PEArray.scala 198:59 PEArray.scala 200:17]
  wire [9:0] _GEN_330 = _T_24 ? 10'h0 : _GEN_127; // @[PEArray.scala 202:32 PEArray.scala 203:15]
  wire [2:0] _GEN_331 = _T_24 ? 3'h0 : state; // @[PEArray.scala 202:32 PEArray.scala 204:15 PEArray.scala 100:22]
  wire [9:0] _GEN_865 = {{4'd0}, GRU_out_width}; // @[PEArray.scala 220:19]
  wire [9:0] _GEN_0 = count % _GEN_865; // @[PEArray.scala 220:19]
  wire [5:0] _T_36 = _GEN_0[5:0]; // @[PEArray.scala 220:19]
  wire [5:0] _T_38 = GRU_out_width - 6'h1; // @[PEArray.scala 220:55]
  wire [5:0] _GEN_334 = _T_36 == _T_38 ? _L0Index_T_2 : 6'h0; // @[PEArray.scala 220:62 PEArray.scala 221:17 PEArray.scala 214:15]
  wire [5:0] _GEN_346 = _T_41 ? _GEN_334 : L0Index; // @[Conditional.scala 39:67 PEArray.scala 39:24]
  wire [9:0] _GEN_347 = _T_41 ? _GEN_330 : count; // @[Conditional.scala 39:67 PEArray.scala 101:22]
  wire [2:0] _GEN_348 = _T_41 ? _GEN_331 : state; // @[Conditional.scala 39:67 PEArray.scala 100:22]
  wire [5:0] _GEN_353 = _T_31 ? _GEN_334 : _GEN_346; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_354 = _T_31 ? _GEN_330 : _GEN_347; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_355 = _T_31 ? _GEN_331 : _GEN_348; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_356 = _T_22 ? _GEN_330 : _GEN_354; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_357 = _T_22 ? _GEN_329 : _GEN_353; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_458 = _T_22 ? _GEN_331 : _GEN_355; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_690 = _T_3 ? _GEN_118 : {{2'd0}, GRU_out_width}; // @[Conditional.scala 40:58 PEArray.scala 104:26]
  FP16MulAdder FP16MAC ( // @[PEArray.scala 72:23]
    .io_a(FP16MAC_io_a),
    .io_b(FP16MAC_io_b),
    .io_c(FP16MAC_io_c),
    .io_out(FP16MAC_io_out)
  );
  assign io_ToBelowPE = mux2out_reg; // @[PEArray.scala 94:16]
  assign FP16MAC_io_a = sel1 ? io_FromL1 : io_FromLeftPE; // @[PEArray.scala 50:14 PEArray.scala 50:23 PEArray.scala 51:24]
  assign FP16MAC_io_b = sel5 ? mux4out : _GEN_105; // @[PEArray.scala 77:13 PEArray.scala 78:18 PEArray.scala 81:18]
  assign FP16MAC_io_c = sel5 ? _GEN_105 : mux4out; // @[PEArray.scala 77:13 PEArray.scala 79:18 PEArray.scala 82:18]
  always @(posedge clock) begin
    if (reset) begin // @[PEArray.scala 39:24]
      L0Index <= 6'h0; // @[PEArray.scala 39:24]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h1; // @[PEArray.scala 159:15]
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        L0Index <= 6'he; // @[PEArray.scala 181:15]
      end else begin
        L0Index <= _GEN_357;
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_0 <= _GEN_229;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_1 <= _GEN_230;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_2 <= _GEN_231;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_3 <= _GEN_232;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_4 <= _GEN_233;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_5 <= _GEN_234;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_6 <= _GEN_235;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_7 <= _GEN_236;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_8 <= _GEN_237;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_9 <= _GEN_238;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_10 <= _GEN_239;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_11 <= _GEN_240;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_12 <= _GEN_241;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_13 <= _GEN_242;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_14 <= _GEN_243;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_15 <= _GEN_244;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_16 <= _GEN_245;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_17 <= _GEN_246;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_18 <= _GEN_247;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_19 <= _GEN_248;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_20 <= _GEN_249;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_21 <= _GEN_250;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_22 <= _GEN_251;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_23 <= _GEN_252;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_24 <= _GEN_253;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_25 <= _GEN_254;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_26 <= _GEN_255;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_27 <= _GEN_256;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_28 <= _GEN_257;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_29 <= _GEN_258;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_30 <= _GEN_259;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_31 <= _GEN_260;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_32 <= _GEN_261;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_33 <= _GEN_262;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_34 <= _GEN_263;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_35 <= _GEN_264;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_36 <= _GEN_265;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_37 <= _GEN_266;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_38 <= _GEN_267;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_39 <= _GEN_268;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_40 <= _GEN_269;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_41 <= _GEN_270;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_42 <= _GEN_271;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_43 <= _GEN_272;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_44 <= _GEN_273;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_45 <= _GEN_274;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_46 <= _GEN_275;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_47 <= _GEN_276;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_48 <= _GEN_277;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_49 <= _GEN_278;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_50 <= _GEN_279;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_51 <= _GEN_280;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_52 <= _GEN_281;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_53 <= _GEN_282;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_54 <= _GEN_283;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_55 <= _GEN_284;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_56 <= _GEN_285;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_57 <= _GEN_286;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_58 <= _GEN_287;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_59 <= _GEN_288;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_60 <= _GEN_289;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_61 <= _GEN_290;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_62 <= _GEN_291;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_63 <= _GEN_292;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_64 <= _GEN_293;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_65 <= _GEN_294;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_66 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_67 <= _GEN_296;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_68 <= _GEN_297;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_69 <= _GEN_298;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_70 <= _GEN_299;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_71 <= _GEN_300;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_72 <= _GEN_301;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_73 <= _GEN_302;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_74 <= _GEN_303;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_75 <= _GEN_304;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_76 <= _GEN_305;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_77 <= _GEN_306;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_78 <= _GEN_307;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_79 <= _GEN_308;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_80 <= _GEN_309;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_81 <= _GEN_310;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_82 <= _GEN_311;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_83 <= _GEN_312;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_84 <= _GEN_313;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_85 <= _GEN_314;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_86 <= _GEN_315;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_87 <= _GEN_316;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_88 <= _GEN_317;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_89 <= _GEN_318;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_90 <= _GEN_319;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_91 <= _GEN_320;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_92 <= _GEN_321;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_93 <= _GEN_322;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_94 <= _GEN_323;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_95 <= _GEN_324;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_96 <= _GEN_325;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_97 <= _GEN_326;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_98 <= _GEN_327;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_99 <= _GEN_328;
          end
        end
      end
    end
    if (reset) begin // @[PEArray.scala 100:22]
      state <= 3'h0; // @[PEArray.scala 100:22]
    end else if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[0]) begin // @[PEArray.scala 116:57]
        state <= 3'h1;
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      if (count == 10'h33) begin // @[PEArray.scala 164:27]
        state <= 3'h0; // @[PEArray.scala 166:15]
      end
    end else if (_T_16) begin // @[Conditional.scala 39:67]
      state <= _GEN_126;
    end else begin
      state <= _GEN_458;
    end
    if (reset) begin // @[PEArray.scala 90:28]
      mux2out_reg <= 16'h0; // @[PEArray.scala 90:28]
    end else begin
      mux2out_reg <= MAC_out; // @[PEArray.scala 90:28]
    end
    if (reset) begin // @[PEArray.scala 101:22]
      count <= 10'h0; // @[PEArray.scala 101:22]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        if (count == 10'h33) begin // @[PEArray.scala 164:27]
          count <= 10'h0; // @[PEArray.scala 165:15]
        end else begin
          count <= _GEN_120;
        end
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        count <= _GEN_125;
      end else begin
        count <= _GEN_356;
      end
    end
    GRU_out_width <= _GEN_690[5:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  L0Index = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  L0Memory_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  L0Memory_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  L0Memory_2 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  L0Memory_3 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  L0Memory_4 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  L0Memory_5 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  L0Memory_6 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  L0Memory_7 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  L0Memory_8 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  L0Memory_9 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  L0Memory_10 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  L0Memory_11 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  L0Memory_12 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  L0Memory_13 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  L0Memory_14 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  L0Memory_15 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  L0Memory_16 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  L0Memory_17 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  L0Memory_18 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  L0Memory_19 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  L0Memory_20 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  L0Memory_21 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  L0Memory_22 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  L0Memory_23 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  L0Memory_24 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  L0Memory_25 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  L0Memory_26 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  L0Memory_27 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  L0Memory_28 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  L0Memory_29 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  L0Memory_30 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  L0Memory_31 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  L0Memory_32 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  L0Memory_33 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  L0Memory_34 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  L0Memory_35 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  L0Memory_36 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  L0Memory_37 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  L0Memory_38 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  L0Memory_39 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  L0Memory_40 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  L0Memory_41 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  L0Memory_42 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  L0Memory_43 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  L0Memory_44 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  L0Memory_45 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  L0Memory_46 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  L0Memory_47 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  L0Memory_48 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  L0Memory_49 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  L0Memory_50 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  L0Memory_51 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  L0Memory_52 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  L0Memory_53 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  L0Memory_54 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  L0Memory_55 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  L0Memory_56 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  L0Memory_57 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  L0Memory_58 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  L0Memory_59 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  L0Memory_60 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  L0Memory_61 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  L0Memory_62 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  L0Memory_63 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  L0Memory_64 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  L0Memory_65 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  L0Memory_66 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  L0Memory_67 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  L0Memory_68 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  L0Memory_69 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  L0Memory_70 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  L0Memory_71 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  L0Memory_72 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  L0Memory_73 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  L0Memory_74 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  L0Memory_75 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  L0Memory_76 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  L0Memory_77 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  L0Memory_78 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  L0Memory_79 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  L0Memory_80 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  L0Memory_81 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  L0Memory_82 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  L0Memory_83 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  L0Memory_84 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  L0Memory_85 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  L0Memory_86 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  L0Memory_87 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  L0Memory_88 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  L0Memory_89 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  L0Memory_90 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  L0Memory_91 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  L0Memory_92 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  L0Memory_93 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  L0Memory_94 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  L0Memory_95 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  L0Memory_96 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  L0Memory_97 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  L0Memory_98 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  L0Memory_99 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  state = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  mux2out_reg = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  count = _RAND_103[9:0];
  _RAND_104 = {1{`RANDOM}};
  GRU_out_width = _RAND_104[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PE_35(
  input         clock,
  input         reset,
  input  [15:0] io_FromAbovePE,
  input  [15:0] io_FromLeftPE,
  input  [15:0] io_FromL1,
  input  [2:0]  io_control_signal_control,
  input  [9:0]  io_control_signal_count,
  input  [5:0]  io_control_signal_L0index,
  input  [11:0] io_control_signal_mask,
  input  [7:0]  io_control_signal_gru_out_width,
  output [15:0] io_ToRightPE,
  output [15:0] io_ToBelowPE
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] FP16MAC_io_a; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_b; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_c; // @[PEArray.scala 72:23]
  wire [15:0] FP16MAC_io_out; // @[PEArray.scala 72:23]
  reg [5:0] L0Index; // @[PEArray.scala 39:24]
  reg [15:0] L0Memory_0; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_1; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_2; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_3; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_4; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_5; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_6; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_7; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_8; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_9; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_10; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_11; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_12; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_13; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_14; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_15; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_16; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_17; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_18; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_19; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_20; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_21; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_22; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_23; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_24; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_25; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_26; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_27; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_28; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_29; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_30; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_31; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_32; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_33; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_34; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_35; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_36; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_37; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_38; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_39; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_40; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_41; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_42; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_43; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_44; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_45; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_46; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_47; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_48; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_49; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_50; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_51; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_52; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_53; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_54; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_55; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_56; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_57; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_58; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_59; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_60; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_61; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_62; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_63; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_64; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_65; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_66; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_67; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_68; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_69; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_70; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_71; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_72; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_73; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_74; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_75; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_76; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_77; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_78; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_79; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_80; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_81; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_82; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_83; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_84; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_85; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_86; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_87; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_88; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_89; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_90; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_91; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_92; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_93; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_94; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_95; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_96; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_97; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_98; // @[PEArray.scala 40:21]
  reg [15:0] L0Memory_99; // @[PEArray.scala 40:21]
  reg [2:0] state; // @[PEArray.scala 100:22]
  wire  _T_3 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_12 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_16 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_22 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_31 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_41 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_342 = _T_41 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 231:12 PEArray.scala 32:8]
  wire  _GEN_349 = _T_31 ? 1'h0 : _GEN_342; // @[Conditional.scala 39:67 PEArray.scala 208:12]
  wire  _GEN_459 = _T_22 | _GEN_349; // @[Conditional.scala 39:67 PEArray.scala 32:8]
  wire  _GEN_463 = _T_16 ? 1'h0 : _GEN_459; // @[Conditional.scala 39:67]
  wire  _GEN_572 = _T_12 | _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 149:12]
  wire  sel1 = _T_3 | _GEN_572; // @[Conditional.scala 40:58 PEArray.scala 108:12]
  wire [15:0] MAC_out = FP16MAC_io_out; // @[PEArray.scala 47:21 PEArray.scala 85:11]
  wire  _GEN_465 = _T_16 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 PEArray.scala 177:12]
  wire  _GEN_580 = _T_12 | _GEN_465; // @[Conditional.scala 39:67 PEArray.scala 34:8]
  wire  sel3 = _T_3 | _GEN_580; // @[Conditional.scala 40:58 PEArray.scala 110:12]
  wire [1:0] _GEN_344 = _T_41 ? 2'h2 : 2'h0; // @[Conditional.scala 39:67 PEArray.scala 233:12 PEArray.scala 35:8]
  wire [1:0] _GEN_351 = _T_31 ? 2'h2 : _GEN_344; // @[Conditional.scala 39:67 PEArray.scala 210:12]
  wire [1:0] _GEN_461 = _T_22 ? 2'h0 : _GEN_351; // @[Conditional.scala 39:67 PEArray.scala 35:8]
  wire [1:0] _GEN_466 = _T_16 ? 2'h0 : _GEN_461; // @[Conditional.scala 39:67 PEArray.scala 178:12]
  wire [1:0] _GEN_574 = _T_12 ? 2'h1 : _GEN_466; // @[Conditional.scala 39:67]
  wire [1:0] sel4 = _T_3 ? 2'h0 : _GEN_574; // @[Conditional.scala 40:58 PEArray.scala 111:12]
  wire [15:0] _GEN_3 = sel4 == 2'h2 ? io_FromL1 : 16'h0; // @[PEArray.scala 65:28 PEArray.scala 66:15 PEArray.scala 69:15]
  wire [15:0] _GEN_4 = sel4 == 2'h1 ? io_FromAbovePE : _GEN_3; // @[PEArray.scala 62:28 PEArray.scala 63:15]
  wire [15:0] mux4out = sel4 == 2'h0 ? 16'h0 : _GEN_4; // @[PEArray.scala 59:22 PEArray.scala 60:13]
  wire [15:0] _GEN_7 = 6'h1 == L0Index ? L0Memory_1 : L0Memory_0; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_8 = 6'h2 == L0Index ? L0Memory_2 : _GEN_7; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_9 = 6'h3 == L0Index ? L0Memory_3 : _GEN_8; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_10 = 6'h4 == L0Index ? L0Memory_4 : _GEN_9; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_11 = 6'h5 == L0Index ? L0Memory_5 : _GEN_10; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_12 = 6'h6 == L0Index ? L0Memory_6 : _GEN_11; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_13 = 6'h7 == L0Index ? L0Memory_7 : _GEN_12; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_14 = 6'h8 == L0Index ? L0Memory_8 : _GEN_13; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_15 = 6'h9 == L0Index ? L0Memory_9 : _GEN_14; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_16 = 6'ha == L0Index ? L0Memory_10 : _GEN_15; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_17 = 6'hb == L0Index ? L0Memory_11 : _GEN_16; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_18 = 6'hc == L0Index ? L0Memory_12 : _GEN_17; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_19 = 6'hd == L0Index ? L0Memory_13 : _GEN_18; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_20 = 6'he == L0Index ? L0Memory_14 : _GEN_19; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_21 = 6'hf == L0Index ? L0Memory_15 : _GEN_20; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_22 = 6'h10 == L0Index ? L0Memory_16 : _GEN_21; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_23 = 6'h11 == L0Index ? L0Memory_17 : _GEN_22; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_24 = 6'h12 == L0Index ? L0Memory_18 : _GEN_23; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_25 = 6'h13 == L0Index ? L0Memory_19 : _GEN_24; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_26 = 6'h14 == L0Index ? L0Memory_20 : _GEN_25; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_27 = 6'h15 == L0Index ? L0Memory_21 : _GEN_26; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_28 = 6'h16 == L0Index ? L0Memory_22 : _GEN_27; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_29 = 6'h17 == L0Index ? L0Memory_23 : _GEN_28; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_30 = 6'h18 == L0Index ? L0Memory_24 : _GEN_29; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_31 = 6'h19 == L0Index ? L0Memory_25 : _GEN_30; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_32 = 6'h1a == L0Index ? L0Memory_26 : _GEN_31; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_33 = 6'h1b == L0Index ? L0Memory_27 : _GEN_32; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_34 = 6'h1c == L0Index ? L0Memory_28 : _GEN_33; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_35 = 6'h1d == L0Index ? L0Memory_29 : _GEN_34; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_36 = 6'h1e == L0Index ? L0Memory_30 : _GEN_35; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_37 = 6'h1f == L0Index ? L0Memory_31 : _GEN_36; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_38 = 6'h20 == L0Index ? L0Memory_32 : _GEN_37; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_39 = 6'h21 == L0Index ? L0Memory_33 : _GEN_38; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_40 = 6'h22 == L0Index ? L0Memory_34 : _GEN_39; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_41 = 6'h23 == L0Index ? L0Memory_35 : _GEN_40; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_42 = 6'h24 == L0Index ? L0Memory_36 : _GEN_41; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_43 = 6'h25 == L0Index ? L0Memory_37 : _GEN_42; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_44 = 6'h26 == L0Index ? L0Memory_38 : _GEN_43; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_45 = 6'h27 == L0Index ? L0Memory_39 : _GEN_44; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_46 = 6'h28 == L0Index ? L0Memory_40 : _GEN_45; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_47 = 6'h29 == L0Index ? L0Memory_41 : _GEN_46; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_48 = 6'h2a == L0Index ? L0Memory_42 : _GEN_47; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_49 = 6'h2b == L0Index ? L0Memory_43 : _GEN_48; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_50 = 6'h2c == L0Index ? L0Memory_44 : _GEN_49; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_51 = 6'h2d == L0Index ? L0Memory_45 : _GEN_50; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_52 = 6'h2e == L0Index ? L0Memory_46 : _GEN_51; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_53 = 6'h2f == L0Index ? L0Memory_47 : _GEN_52; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_54 = 6'h30 == L0Index ? L0Memory_48 : _GEN_53; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_55 = 6'h31 == L0Index ? L0Memory_49 : _GEN_54; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_56 = 6'h32 == L0Index ? L0Memory_50 : _GEN_55; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_57 = 6'h33 == L0Index ? L0Memory_51 : _GEN_56; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_58 = 6'h34 == L0Index ? L0Memory_52 : _GEN_57; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_59 = 6'h35 == L0Index ? L0Memory_53 : _GEN_58; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_60 = 6'h36 == L0Index ? L0Memory_54 : _GEN_59; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_61 = 6'h37 == L0Index ? L0Memory_55 : _GEN_60; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_62 = 6'h38 == L0Index ? L0Memory_56 : _GEN_61; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_63 = 6'h39 == L0Index ? L0Memory_57 : _GEN_62; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_64 = 6'h3a == L0Index ? L0Memory_58 : _GEN_63; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_65 = 6'h3b == L0Index ? L0Memory_59 : _GEN_64; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_66 = 6'h3c == L0Index ? L0Memory_60 : _GEN_65; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_67 = 6'h3d == L0Index ? L0Memory_61 : _GEN_66; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_68 = 6'h3e == L0Index ? L0Memory_62 : _GEN_67; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_69 = 6'h3f == L0Index ? L0Memory_63 : _GEN_68; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [6:0] _GEN_793 = {{1'd0}, L0Index}; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_70 = 7'h40 == _GEN_793 ? L0Memory_64 : _GEN_69; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_71 = 7'h41 == _GEN_793 ? L0Memory_65 : _GEN_70; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_72 = 7'h42 == _GEN_793 ? L0Memory_66 : _GEN_71; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_73 = 7'h43 == _GEN_793 ? L0Memory_67 : _GEN_72; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_74 = 7'h44 == _GEN_793 ? L0Memory_68 : _GEN_73; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_75 = 7'h45 == _GEN_793 ? L0Memory_69 : _GEN_74; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_76 = 7'h46 == _GEN_793 ? L0Memory_70 : _GEN_75; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_77 = 7'h47 == _GEN_793 ? L0Memory_71 : _GEN_76; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_78 = 7'h48 == _GEN_793 ? L0Memory_72 : _GEN_77; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_79 = 7'h49 == _GEN_793 ? L0Memory_73 : _GEN_78; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_80 = 7'h4a == _GEN_793 ? L0Memory_74 : _GEN_79; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_81 = 7'h4b == _GEN_793 ? L0Memory_75 : _GEN_80; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_82 = 7'h4c == _GEN_793 ? L0Memory_76 : _GEN_81; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_83 = 7'h4d == _GEN_793 ? L0Memory_77 : _GEN_82; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_84 = 7'h4e == _GEN_793 ? L0Memory_78 : _GEN_83; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_85 = 7'h4f == _GEN_793 ? L0Memory_79 : _GEN_84; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_86 = 7'h50 == _GEN_793 ? L0Memory_80 : _GEN_85; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_87 = 7'h51 == _GEN_793 ? L0Memory_81 : _GEN_86; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_88 = 7'h52 == _GEN_793 ? L0Memory_82 : _GEN_87; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_89 = 7'h53 == _GEN_793 ? L0Memory_83 : _GEN_88; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_90 = 7'h54 == _GEN_793 ? L0Memory_84 : _GEN_89; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_91 = 7'h55 == _GEN_793 ? L0Memory_85 : _GEN_90; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_92 = 7'h56 == _GEN_793 ? L0Memory_86 : _GEN_91; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_93 = 7'h57 == _GEN_793 ? L0Memory_87 : _GEN_92; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_94 = 7'h58 == _GEN_793 ? L0Memory_88 : _GEN_93; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_95 = 7'h59 == _GEN_793 ? L0Memory_89 : _GEN_94; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_96 = 7'h5a == _GEN_793 ? L0Memory_90 : _GEN_95; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_97 = 7'h5b == _GEN_793 ? L0Memory_91 : _GEN_96; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_98 = 7'h5c == _GEN_793 ? L0Memory_92 : _GEN_97; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_99 = 7'h5d == _GEN_793 ? L0Memory_93 : _GEN_98; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_100 = 7'h5e == _GEN_793 ? L0Memory_94 : _GEN_99; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_101 = 7'h5f == _GEN_793 ? L0Memory_95 : _GEN_100; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_102 = 7'h60 == _GEN_793 ? L0Memory_96 : _GEN_101; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_103 = 7'h61 == _GEN_793 ? L0Memory_97 : _GEN_102; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_104 = 7'h62 == _GEN_793 ? L0Memory_98 : _GEN_103; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire [15:0] _GEN_105 = 7'h63 == _GEN_793 ? L0Memory_99 : _GEN_104; // @[PEArray.scala 79:18 PEArray.scala 79:18]
  wire  _GEN_575 = _T_12 ? 1'h0 : _GEN_463; // @[Conditional.scala 39:67 PEArray.scala 157:12]
  wire  sel5 = _T_3 ? 1'h0 : _GEN_575; // @[Conditional.scala 40:58 PEArray.scala 112:12]
  reg [15:0] mux2out_reg; // @[PEArray.scala 90:28]
  reg [15:0] mux3out_reg; // @[PEArray.scala 91:28]
  reg [9:0] count; // @[PEArray.scala 101:22]
  reg [9:0] count_max; // @[PEArray.scala 102:22]
  reg [5:0] L0index_begin; // @[PEArray.scala 103:26]
  reg [5:0] GRU_out_width; // @[PEArray.scala 104:26]
  wire  _T_6 = 3'h0 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_7 = 3'h1 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_8 = 3'h2 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_9 = 3'h3 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_10 = 3'h4 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire  _T_11 = 3'h5 == io_control_signal_control; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_109 = _T_11 ? 3'h5 : state; // @[Conditional.scala 39:67 PEArray.scala 140:19 PEArray.scala 100:22]
  wire [2:0] _GEN_110 = _T_10 ? 3'h4 : _GEN_109; // @[Conditional.scala 39:67 PEArray.scala 136:19]
  wire [2:0] _GEN_111 = _T_9 ? 3'h3 : _GEN_110; // @[Conditional.scala 39:67 PEArray.scala 132:19]
  wire [2:0] _GEN_112 = _T_8 ? 3'h2 : _GEN_111; // @[Conditional.scala 39:67 PEArray.scala 128:19]
  wire [2:0] _GEN_113 = _T_7 ? 3'h1 : _GEN_112; // @[Conditional.scala 39:67 PEArray.scala 124:19]
  wire [7:0] _GEN_118 = io_control_signal_mask[0] ? io_control_signal_gru_out_width : {{2'd0}, GRU_out_width}; // @[PEArray.scala 116:57 PEArray.scala 145:23 PEArray.scala 104:26]
  wire [9:0] _count_T_1 = count + 10'h1; // @[PEArray.scala 162:24]
  wire [9:0] _GEN_120 = count != 10'h33 ? _count_T_1 : count; // @[PEArray.scala 161:27 PEArray.scala 162:15 PEArray.scala 101:22]
  wire [9:0] _GEN_124 = count != 10'h188 ? _count_T_1 : count; // @[PEArray.scala 183:28 PEArray.scala 184:15 PEArray.scala 101:22]
  wire [9:0] _GEN_125 = count == 10'h188 ? 10'h0 : _GEN_124; // @[PEArray.scala 186:28 PEArray.scala 187:15]
  wire [2:0] _GEN_126 = count == 10'h188 ? 3'h0 : state; // @[PEArray.scala 186:28 PEArray.scala 188:15 PEArray.scala 100:22]
  wire [9:0] _GEN_127 = count != count_max ? _count_T_1 : count; // @[PEArray.scala 192:32 PEArray.scala 193:15 PEArray.scala 101:22]
  wire [5:0] _GEN_128 = count == 10'h0 ? L0index_begin : L0Index; // @[PEArray.scala 195:26 PEArray.scala 196:17 PEArray.scala 39:24]
  wire [9:0] _T_27 = count_max - 10'h1; // @[PEArray.scala 198:51]
  wire [15:0] _GEN_129 = 6'h0 == L0Index ? io_FromL1 : L0Memory_0; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_130 = 6'h1 == L0Index ? io_FromL1 : L0Memory_1; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_131 = 6'h2 == L0Index ? io_FromL1 : L0Memory_2; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_132 = 6'h3 == L0Index ? io_FromL1 : L0Memory_3; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_133 = 6'h4 == L0Index ? io_FromL1 : L0Memory_4; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_134 = 6'h5 == L0Index ? io_FromL1 : L0Memory_5; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_135 = 6'h6 == L0Index ? io_FromL1 : L0Memory_6; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_136 = 6'h7 == L0Index ? io_FromL1 : L0Memory_7; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_137 = 6'h8 == L0Index ? io_FromL1 : L0Memory_8; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_138 = 6'h9 == L0Index ? io_FromL1 : L0Memory_9; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_139 = 6'ha == L0Index ? io_FromL1 : L0Memory_10; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_140 = 6'hb == L0Index ? io_FromL1 : L0Memory_11; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_141 = 6'hc == L0Index ? io_FromL1 : L0Memory_12; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_142 = 6'hd == L0Index ? io_FromL1 : L0Memory_13; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_143 = 6'he == L0Index ? io_FromL1 : L0Memory_14; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_144 = 6'hf == L0Index ? io_FromL1 : L0Memory_15; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_145 = 6'h10 == L0Index ? io_FromL1 : L0Memory_16; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_146 = 6'h11 == L0Index ? io_FromL1 : L0Memory_17; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_147 = 6'h12 == L0Index ? io_FromL1 : L0Memory_18; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_148 = 6'h13 == L0Index ? io_FromL1 : L0Memory_19; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_149 = 6'h14 == L0Index ? io_FromL1 : L0Memory_20; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_150 = 6'h15 == L0Index ? io_FromL1 : L0Memory_21; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_151 = 6'h16 == L0Index ? io_FromL1 : L0Memory_22; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_152 = 6'h17 == L0Index ? io_FromL1 : L0Memory_23; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_153 = 6'h18 == L0Index ? io_FromL1 : L0Memory_24; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_154 = 6'h19 == L0Index ? io_FromL1 : L0Memory_25; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_155 = 6'h1a == L0Index ? io_FromL1 : L0Memory_26; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_156 = 6'h1b == L0Index ? io_FromL1 : L0Memory_27; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_157 = 6'h1c == L0Index ? io_FromL1 : L0Memory_28; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_158 = 6'h1d == L0Index ? io_FromL1 : L0Memory_29; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_159 = 6'h1e == L0Index ? io_FromL1 : L0Memory_30; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_160 = 6'h1f == L0Index ? io_FromL1 : L0Memory_31; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_161 = 6'h20 == L0Index ? io_FromL1 : L0Memory_32; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_162 = 6'h21 == L0Index ? io_FromL1 : L0Memory_33; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_163 = 6'h22 == L0Index ? io_FromL1 : L0Memory_34; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_164 = 6'h23 == L0Index ? io_FromL1 : L0Memory_35; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_165 = 6'h24 == L0Index ? io_FromL1 : L0Memory_36; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_166 = 6'h25 == L0Index ? io_FromL1 : L0Memory_37; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_167 = 6'h26 == L0Index ? io_FromL1 : L0Memory_38; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_168 = 6'h27 == L0Index ? io_FromL1 : L0Memory_39; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_169 = 6'h28 == L0Index ? io_FromL1 : L0Memory_40; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_170 = 6'h29 == L0Index ? io_FromL1 : L0Memory_41; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_171 = 6'h2a == L0Index ? io_FromL1 : L0Memory_42; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_172 = 6'h2b == L0Index ? io_FromL1 : L0Memory_43; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_173 = 6'h2c == L0Index ? io_FromL1 : L0Memory_44; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_174 = 6'h2d == L0Index ? io_FromL1 : L0Memory_45; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_175 = 6'h2e == L0Index ? io_FromL1 : L0Memory_46; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_176 = 6'h2f == L0Index ? io_FromL1 : L0Memory_47; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_177 = 6'h30 == L0Index ? io_FromL1 : L0Memory_48; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_178 = 6'h31 == L0Index ? io_FromL1 : L0Memory_49; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_179 = 6'h32 == L0Index ? io_FromL1 : L0Memory_50; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_180 = 6'h33 == L0Index ? io_FromL1 : L0Memory_51; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_181 = 6'h34 == L0Index ? io_FromL1 : L0Memory_52; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_182 = 6'h35 == L0Index ? io_FromL1 : L0Memory_53; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_183 = 6'h36 == L0Index ? io_FromL1 : L0Memory_54; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_184 = 6'h37 == L0Index ? io_FromL1 : L0Memory_55; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_185 = 6'h38 == L0Index ? io_FromL1 : L0Memory_56; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_186 = 6'h39 == L0Index ? io_FromL1 : L0Memory_57; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_187 = 6'h3a == L0Index ? io_FromL1 : L0Memory_58; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_188 = 6'h3b == L0Index ? io_FromL1 : L0Memory_59; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_189 = 6'h3c == L0Index ? io_FromL1 : L0Memory_60; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_190 = 6'h3d == L0Index ? io_FromL1 : L0Memory_61; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_191 = 6'h3e == L0Index ? io_FromL1 : L0Memory_62; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_192 = 6'h3f == L0Index ? io_FromL1 : L0Memory_63; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_193 = 7'h40 == _GEN_793 ? io_FromL1 : L0Memory_64; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_194 = 7'h41 == _GEN_793 ? io_FromL1 : L0Memory_65; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_195 = 7'h42 == _GEN_793 ? io_FromL1 : L0Memory_66; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_196 = 7'h43 == _GEN_793 ? io_FromL1 : L0Memory_67; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_197 = 7'h44 == _GEN_793 ? io_FromL1 : L0Memory_68; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_198 = 7'h45 == _GEN_793 ? io_FromL1 : L0Memory_69; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_199 = 7'h46 == _GEN_793 ? io_FromL1 : L0Memory_70; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_200 = 7'h47 == _GEN_793 ? io_FromL1 : L0Memory_71; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_201 = 7'h48 == _GEN_793 ? io_FromL1 : L0Memory_72; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_202 = 7'h49 == _GEN_793 ? io_FromL1 : L0Memory_73; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_203 = 7'h4a == _GEN_793 ? io_FromL1 : L0Memory_74; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_204 = 7'h4b == _GEN_793 ? io_FromL1 : L0Memory_75; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_205 = 7'h4c == _GEN_793 ? io_FromL1 : L0Memory_76; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_206 = 7'h4d == _GEN_793 ? io_FromL1 : L0Memory_77; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_207 = 7'h4e == _GEN_793 ? io_FromL1 : L0Memory_78; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_208 = 7'h4f == _GEN_793 ? io_FromL1 : L0Memory_79; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_209 = 7'h50 == _GEN_793 ? io_FromL1 : L0Memory_80; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_210 = 7'h51 == _GEN_793 ? io_FromL1 : L0Memory_81; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_211 = 7'h52 == _GEN_793 ? io_FromL1 : L0Memory_82; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_212 = 7'h53 == _GEN_793 ? io_FromL1 : L0Memory_83; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_213 = 7'h54 == _GEN_793 ? io_FromL1 : L0Memory_84; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_214 = 7'h55 == _GEN_793 ? io_FromL1 : L0Memory_85; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_215 = 7'h56 == _GEN_793 ? io_FromL1 : L0Memory_86; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_216 = 7'h57 == _GEN_793 ? io_FromL1 : L0Memory_87; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_217 = 7'h58 == _GEN_793 ? io_FromL1 : L0Memory_88; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_218 = 7'h59 == _GEN_793 ? io_FromL1 : L0Memory_89; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_219 = 7'h5a == _GEN_793 ? io_FromL1 : L0Memory_90; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_220 = 7'h5b == _GEN_793 ? io_FromL1 : L0Memory_91; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_221 = 7'h5c == _GEN_793 ? io_FromL1 : L0Memory_92; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_222 = 7'h5d == _GEN_793 ? io_FromL1 : L0Memory_93; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_223 = 7'h5e == _GEN_793 ? io_FromL1 : L0Memory_94; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_224 = 7'h5f == _GEN_793 ? io_FromL1 : L0Memory_95; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_225 = 7'h60 == _GEN_793 ? io_FromL1 : L0Memory_96; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_226 = 7'h61 == _GEN_793 ? io_FromL1 : L0Memory_97; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_227 = 7'h62 == _GEN_793 ? io_FromL1 : L0Memory_98; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [15:0] _GEN_228 = 7'h63 == _GEN_793 ? io_FromL1 : L0Memory_99; // @[PEArray.scala 199:27 PEArray.scala 199:27 PEArray.scala 40:21]
  wire [5:0] _L0Index_T_2 = L0Index + 6'h1; // @[PEArray.scala 200:28]
  wire [15:0] _GEN_229 = count >= 10'h1 & count <= _T_27 ? _GEN_129 : L0Memory_0; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_230 = count >= 10'h1 & count <= _T_27 ? _GEN_130 : L0Memory_1; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_231 = count >= 10'h1 & count <= _T_27 ? _GEN_131 : L0Memory_2; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_232 = count >= 10'h1 & count <= _T_27 ? _GEN_132 : L0Memory_3; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_233 = count >= 10'h1 & count <= _T_27 ? _GEN_133 : L0Memory_4; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_234 = count >= 10'h1 & count <= _T_27 ? _GEN_134 : L0Memory_5; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_235 = count >= 10'h1 & count <= _T_27 ? _GEN_135 : L0Memory_6; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_236 = count >= 10'h1 & count <= _T_27 ? _GEN_136 : L0Memory_7; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_237 = count >= 10'h1 & count <= _T_27 ? _GEN_137 : L0Memory_8; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_238 = count >= 10'h1 & count <= _T_27 ? _GEN_138 : L0Memory_9; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_239 = count >= 10'h1 & count <= _T_27 ? _GEN_139 : L0Memory_10; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_240 = count >= 10'h1 & count <= _T_27 ? _GEN_140 : L0Memory_11; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_241 = count >= 10'h1 & count <= _T_27 ? _GEN_141 : L0Memory_12; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_242 = count >= 10'h1 & count <= _T_27 ? _GEN_142 : L0Memory_13; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_243 = count >= 10'h1 & count <= _T_27 ? _GEN_143 : L0Memory_14; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_244 = count >= 10'h1 & count <= _T_27 ? _GEN_144 : L0Memory_15; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_245 = count >= 10'h1 & count <= _T_27 ? _GEN_145 : L0Memory_16; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_246 = count >= 10'h1 & count <= _T_27 ? _GEN_146 : L0Memory_17; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_247 = count >= 10'h1 & count <= _T_27 ? _GEN_147 : L0Memory_18; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_248 = count >= 10'h1 & count <= _T_27 ? _GEN_148 : L0Memory_19; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_249 = count >= 10'h1 & count <= _T_27 ? _GEN_149 : L0Memory_20; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_250 = count >= 10'h1 & count <= _T_27 ? _GEN_150 : L0Memory_21; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_251 = count >= 10'h1 & count <= _T_27 ? _GEN_151 : L0Memory_22; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_252 = count >= 10'h1 & count <= _T_27 ? _GEN_152 : L0Memory_23; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_253 = count >= 10'h1 & count <= _T_27 ? _GEN_153 : L0Memory_24; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_254 = count >= 10'h1 & count <= _T_27 ? _GEN_154 : L0Memory_25; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_255 = count >= 10'h1 & count <= _T_27 ? _GEN_155 : L0Memory_26; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_256 = count >= 10'h1 & count <= _T_27 ? _GEN_156 : L0Memory_27; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_257 = count >= 10'h1 & count <= _T_27 ? _GEN_157 : L0Memory_28; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_258 = count >= 10'h1 & count <= _T_27 ? _GEN_158 : L0Memory_29; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_259 = count >= 10'h1 & count <= _T_27 ? _GEN_159 : L0Memory_30; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_260 = count >= 10'h1 & count <= _T_27 ? _GEN_160 : L0Memory_31; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_261 = count >= 10'h1 & count <= _T_27 ? _GEN_161 : L0Memory_32; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_262 = count >= 10'h1 & count <= _T_27 ? _GEN_162 : L0Memory_33; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_263 = count >= 10'h1 & count <= _T_27 ? _GEN_163 : L0Memory_34; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_264 = count >= 10'h1 & count <= _T_27 ? _GEN_164 : L0Memory_35; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_265 = count >= 10'h1 & count <= _T_27 ? _GEN_165 : L0Memory_36; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_266 = count >= 10'h1 & count <= _T_27 ? _GEN_166 : L0Memory_37; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_267 = count >= 10'h1 & count <= _T_27 ? _GEN_167 : L0Memory_38; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_268 = count >= 10'h1 & count <= _T_27 ? _GEN_168 : L0Memory_39; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_269 = count >= 10'h1 & count <= _T_27 ? _GEN_169 : L0Memory_40; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_270 = count >= 10'h1 & count <= _T_27 ? _GEN_170 : L0Memory_41; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_271 = count >= 10'h1 & count <= _T_27 ? _GEN_171 : L0Memory_42; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_272 = count >= 10'h1 & count <= _T_27 ? _GEN_172 : L0Memory_43; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_273 = count >= 10'h1 & count <= _T_27 ? _GEN_173 : L0Memory_44; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_274 = count >= 10'h1 & count <= _T_27 ? _GEN_174 : L0Memory_45; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_275 = count >= 10'h1 & count <= _T_27 ? _GEN_175 : L0Memory_46; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_276 = count >= 10'h1 & count <= _T_27 ? _GEN_176 : L0Memory_47; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_277 = count >= 10'h1 & count <= _T_27 ? _GEN_177 : L0Memory_48; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_278 = count >= 10'h1 & count <= _T_27 ? _GEN_178 : L0Memory_49; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_279 = count >= 10'h1 & count <= _T_27 ? _GEN_179 : L0Memory_50; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_280 = count >= 10'h1 & count <= _T_27 ? _GEN_180 : L0Memory_51; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_281 = count >= 10'h1 & count <= _T_27 ? _GEN_181 : L0Memory_52; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_282 = count >= 10'h1 & count <= _T_27 ? _GEN_182 : L0Memory_53; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_283 = count >= 10'h1 & count <= _T_27 ? _GEN_183 : L0Memory_54; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_284 = count >= 10'h1 & count <= _T_27 ? _GEN_184 : L0Memory_55; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_285 = count >= 10'h1 & count <= _T_27 ? _GEN_185 : L0Memory_56; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_286 = count >= 10'h1 & count <= _T_27 ? _GEN_186 : L0Memory_57; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_287 = count >= 10'h1 & count <= _T_27 ? _GEN_187 : L0Memory_58; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_288 = count >= 10'h1 & count <= _T_27 ? _GEN_188 : L0Memory_59; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_289 = count >= 10'h1 & count <= _T_27 ? _GEN_189 : L0Memory_60; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_290 = count >= 10'h1 & count <= _T_27 ? _GEN_190 : L0Memory_61; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_291 = count >= 10'h1 & count <= _T_27 ? _GEN_191 : L0Memory_62; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_292 = count >= 10'h1 & count <= _T_27 ? _GEN_192 : L0Memory_63; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_293 = count >= 10'h1 & count <= _T_27 ? _GEN_193 : L0Memory_64; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_294 = count >= 10'h1 & count <= _T_27 ? _GEN_194 : L0Memory_65; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_295 = count >= 10'h1 & count <= _T_27 ? _GEN_195 : L0Memory_66; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_296 = count >= 10'h1 & count <= _T_27 ? _GEN_196 : L0Memory_67; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_297 = count >= 10'h1 & count <= _T_27 ? _GEN_197 : L0Memory_68; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_298 = count >= 10'h1 & count <= _T_27 ? _GEN_198 : L0Memory_69; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_299 = count >= 10'h1 & count <= _T_27 ? _GEN_199 : L0Memory_70; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_300 = count >= 10'h1 & count <= _T_27 ? _GEN_200 : L0Memory_71; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_301 = count >= 10'h1 & count <= _T_27 ? _GEN_201 : L0Memory_72; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_302 = count >= 10'h1 & count <= _T_27 ? _GEN_202 : L0Memory_73; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_303 = count >= 10'h1 & count <= _T_27 ? _GEN_203 : L0Memory_74; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_304 = count >= 10'h1 & count <= _T_27 ? _GEN_204 : L0Memory_75; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_305 = count >= 10'h1 & count <= _T_27 ? _GEN_205 : L0Memory_76; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_306 = count >= 10'h1 & count <= _T_27 ? _GEN_206 : L0Memory_77; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_307 = count >= 10'h1 & count <= _T_27 ? _GEN_207 : L0Memory_78; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_308 = count >= 10'h1 & count <= _T_27 ? _GEN_208 : L0Memory_79; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_309 = count >= 10'h1 & count <= _T_27 ? _GEN_209 : L0Memory_80; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_310 = count >= 10'h1 & count <= _T_27 ? _GEN_210 : L0Memory_81; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_311 = count >= 10'h1 & count <= _T_27 ? _GEN_211 : L0Memory_82; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_312 = count >= 10'h1 & count <= _T_27 ? _GEN_212 : L0Memory_83; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_313 = count >= 10'h1 & count <= _T_27 ? _GEN_213 : L0Memory_84; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_314 = count >= 10'h1 & count <= _T_27 ? _GEN_214 : L0Memory_85; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_315 = count >= 10'h1 & count <= _T_27 ? _GEN_215 : L0Memory_86; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_316 = count >= 10'h1 & count <= _T_27 ? _GEN_216 : L0Memory_87; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_317 = count >= 10'h1 & count <= _T_27 ? _GEN_217 : L0Memory_88; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_318 = count >= 10'h1 & count <= _T_27 ? _GEN_218 : L0Memory_89; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_319 = count >= 10'h1 & count <= _T_27 ? _GEN_219 : L0Memory_90; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_320 = count >= 10'h1 & count <= _T_27 ? _GEN_220 : L0Memory_91; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_321 = count >= 10'h1 & count <= _T_27 ? _GEN_221 : L0Memory_92; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_322 = count >= 10'h1 & count <= _T_27 ? _GEN_222 : L0Memory_93; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_323 = count >= 10'h1 & count <= _T_27 ? _GEN_223 : L0Memory_94; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_324 = count >= 10'h1 & count <= _T_27 ? _GEN_224 : L0Memory_95; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_325 = count >= 10'h1 & count <= _T_27 ? _GEN_225 : L0Memory_96; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_326 = count >= 10'h1 & count <= _T_27 ? _GEN_226 : L0Memory_97; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_327 = count >= 10'h1 & count <= _T_27 ? _GEN_227 : L0Memory_98; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [15:0] _GEN_328 = count >= 10'h1 & count <= _T_27 ? _GEN_228 : L0Memory_99; // @[PEArray.scala 198:59 PEArray.scala 40:21]
  wire [5:0] _GEN_329 = count >= 10'h1 & count <= _T_27 ? _L0Index_T_2 : _GEN_128; // @[PEArray.scala 198:59 PEArray.scala 200:17]
  wire [9:0] _GEN_330 = count == count_max ? 10'h0 : _GEN_127; // @[PEArray.scala 202:32 PEArray.scala 203:15]
  wire [2:0] _GEN_331 = count == count_max ? 3'h0 : state; // @[PEArray.scala 202:32 PEArray.scala 204:15 PEArray.scala 100:22]
  wire [9:0] _GEN_865 = {{4'd0}, GRU_out_width}; // @[PEArray.scala 220:19]
  wire [9:0] _GEN_0 = count % _GEN_865; // @[PEArray.scala 220:19]
  wire [5:0] _T_36 = _GEN_0[5:0]; // @[PEArray.scala 220:19]
  wire [5:0] _T_38 = GRU_out_width - 6'h1; // @[PEArray.scala 220:55]
  wire [5:0] _GEN_334 = _T_36 == _T_38 ? _L0Index_T_2 : L0index_begin; // @[PEArray.scala 220:62 PEArray.scala 221:17 PEArray.scala 214:15]
  wire [5:0] _GEN_346 = _T_41 ? _GEN_334 : L0Index; // @[Conditional.scala 39:67 PEArray.scala 39:24]
  wire [9:0] _GEN_347 = _T_41 ? _GEN_330 : count; // @[Conditional.scala 39:67 PEArray.scala 101:22]
  wire [2:0] _GEN_348 = _T_41 ? _GEN_331 : state; // @[Conditional.scala 39:67 PEArray.scala 100:22]
  wire [5:0] _GEN_353 = _T_31 ? _GEN_334 : _GEN_346; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_354 = _T_31 ? _GEN_330 : _GEN_347; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_355 = _T_31 ? _GEN_331 : _GEN_348; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_356 = _T_22 ? _GEN_330 : _GEN_354; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_357 = _T_22 ? _GEN_329 : _GEN_353; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_458 = _T_22 ? _GEN_331 : _GEN_355; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_690 = _T_3 ? _GEN_118 : {{2'd0}, GRU_out_width}; // @[Conditional.scala 40:58 PEArray.scala 104:26]
  FP16MulAdder FP16MAC ( // @[PEArray.scala 72:23]
    .io_a(FP16MAC_io_a),
    .io_b(FP16MAC_io_b),
    .io_c(FP16MAC_io_c),
    .io_out(FP16MAC_io_out)
  );
  assign io_ToRightPE = mux3out_reg; // @[PEArray.scala 95:16]
  assign io_ToBelowPE = mux2out_reg; // @[PEArray.scala 94:16]
  assign FP16MAC_io_a = sel1 ? io_FromL1 : io_FromLeftPE; // @[PEArray.scala 50:14 PEArray.scala 50:23 PEArray.scala 51:24]
  assign FP16MAC_io_b = sel5 ? mux4out : _GEN_105; // @[PEArray.scala 77:13 PEArray.scala 78:18 PEArray.scala 81:18]
  assign FP16MAC_io_c = sel5 ? _GEN_105 : mux4out; // @[PEArray.scala 77:13 PEArray.scala 79:18 PEArray.scala 82:18]
  always @(posedge clock) begin
    if (reset) begin // @[PEArray.scala 39:24]
      L0Index <= 6'h0; // @[PEArray.scala 39:24]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        L0Index <= 6'h2; // @[PEArray.scala 159:15]
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        L0Index <= 6'he; // @[PEArray.scala 181:15]
      end else begin
        L0Index <= _GEN_357;
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_0 <= _GEN_229;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_1 <= _GEN_230;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_2 <= _GEN_231;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_3 <= _GEN_232;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_4 <= _GEN_233;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_5 <= _GEN_234;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_6 <= _GEN_235;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_7 <= _GEN_236;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_8 <= _GEN_237;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_9 <= _GEN_238;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_10 <= _GEN_239;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_11 <= _GEN_240;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_12 <= _GEN_241;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_13 <= _GEN_242;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_14 <= _GEN_243;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_15 <= _GEN_244;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_16 <= _GEN_245;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_17 <= _GEN_246;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_18 <= _GEN_247;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_19 <= _GEN_248;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_20 <= _GEN_249;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_21 <= _GEN_250;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_22 <= _GEN_251;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_23 <= _GEN_252;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_24 <= _GEN_253;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_25 <= _GEN_254;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_26 <= _GEN_255;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_27 <= _GEN_256;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_28 <= _GEN_257;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_29 <= _GEN_258;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_30 <= _GEN_259;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_31 <= _GEN_260;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_32 <= _GEN_261;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_33 <= _GEN_262;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_34 <= _GEN_263;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_35 <= _GEN_264;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_36 <= _GEN_265;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_37 <= _GEN_266;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_38 <= _GEN_267;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_39 <= _GEN_268;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_40 <= _GEN_269;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_41 <= _GEN_270;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_42 <= _GEN_271;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_43 <= _GEN_272;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_44 <= _GEN_273;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_45 <= _GEN_274;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_46 <= _GEN_275;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_47 <= _GEN_276;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_48 <= _GEN_277;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_49 <= _GEN_278;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_50 <= _GEN_279;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_51 <= _GEN_280;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_52 <= _GEN_281;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_53 <= _GEN_282;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_54 <= _GEN_283;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_55 <= _GEN_284;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_56 <= _GEN_285;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_57 <= _GEN_286;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_58 <= _GEN_287;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_59 <= _GEN_288;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_60 <= _GEN_289;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_61 <= _GEN_290;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_62 <= _GEN_291;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_63 <= _GEN_292;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_64 <= _GEN_293;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_65 <= _GEN_294;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_66 <= _GEN_295;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_67 <= _GEN_296;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_68 <= _GEN_297;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_69 <= _GEN_298;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_70 <= _GEN_299;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_71 <= _GEN_300;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_72 <= _GEN_301;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_73 <= _GEN_302;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_74 <= _GEN_303;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_75 <= _GEN_304;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_76 <= _GEN_305;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_77 <= _GEN_306;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_78 <= _GEN_307;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_79 <= _GEN_308;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_80 <= _GEN_309;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_81 <= _GEN_310;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_82 <= _GEN_311;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_83 <= _GEN_312;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_84 <= _GEN_313;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_85 <= _GEN_314;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_86 <= _GEN_315;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_87 <= _GEN_316;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_88 <= _GEN_317;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_89 <= _GEN_318;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_90 <= _GEN_319;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_91 <= _GEN_320;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_92 <= _GEN_321;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_93 <= _GEN_322;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_94 <= _GEN_323;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_95 <= _GEN_324;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_96 <= _GEN_325;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_97 <= _GEN_326;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_98 <= _GEN_327;
          end
        end
      end
    end
    if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (!(_T_16)) begin // @[Conditional.scala 39:67]
          if (_T_22) begin // @[Conditional.scala 39:67]
            L0Memory_99 <= _GEN_328;
          end
        end
      end
    end
    if (reset) begin // @[PEArray.scala 100:22]
      state <= 3'h0; // @[PEArray.scala 100:22]
    end else if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[0]) begin // @[PEArray.scala 116:57]
        if (_T_6) begin // @[Conditional.scala 40:58]
          state <= 3'h0; // @[PEArray.scala 120:19]
        end else begin
          state <= _GEN_113;
        end
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      if (count == 10'h33) begin // @[PEArray.scala 164:27]
        state <= 3'h0; // @[PEArray.scala 166:15]
      end
    end else if (_T_16) begin // @[Conditional.scala 39:67]
      state <= _GEN_126;
    end else begin
      state <= _GEN_458;
    end
    if (reset) begin // @[PEArray.scala 90:28]
      mux2out_reg <= 16'h0; // @[PEArray.scala 90:28]
    end else begin
      mux2out_reg <= MAC_out; // @[PEArray.scala 90:28]
    end
    if (reset) begin // @[PEArray.scala 91:28]
      mux3out_reg <= 16'h0; // @[PEArray.scala 91:28]
    end else if (sel3) begin // @[PEArray.scala 56:14]
      mux3out_reg <= MAC_out; // @[PEArray.scala 56:23]
    end else if (sel1) begin // @[PEArray.scala 50:14]
      mux3out_reg <= io_FromL1; // @[PEArray.scala 50:23]
    end else begin
      mux3out_reg <= io_FromLeftPE; // @[PEArray.scala 51:24]
    end
    if (reset) begin // @[PEArray.scala 101:22]
      count <= 10'h0; // @[PEArray.scala 101:22]
    end else if (!(_T_3)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        if (count == 10'h33) begin // @[PEArray.scala 164:27]
          count <= 10'h0; // @[PEArray.scala 165:15]
        end else begin
          count <= _GEN_120;
        end
      end else if (_T_16) begin // @[Conditional.scala 39:67]
        count <= _GEN_125;
      end else begin
        count <= _GEN_356;
      end
    end
    if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[0]) begin // @[PEArray.scala 116:57]
        count_max <= io_control_signal_count; // @[PEArray.scala 143:19]
      end
    end
    if (_T_3) begin // @[Conditional.scala 40:58]
      if (io_control_signal_mask[0]) begin // @[PEArray.scala 116:57]
        L0index_begin <= io_control_signal_L0index; // @[PEArray.scala 144:23]
      end
    end
    GRU_out_width <= _GEN_690[5:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  L0Index = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  L0Memory_0 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  L0Memory_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  L0Memory_2 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  L0Memory_3 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  L0Memory_4 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  L0Memory_5 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  L0Memory_6 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  L0Memory_7 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  L0Memory_8 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  L0Memory_9 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  L0Memory_10 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  L0Memory_11 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  L0Memory_12 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  L0Memory_13 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  L0Memory_14 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  L0Memory_15 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  L0Memory_16 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  L0Memory_17 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  L0Memory_18 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  L0Memory_19 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  L0Memory_20 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  L0Memory_21 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  L0Memory_22 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  L0Memory_23 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  L0Memory_24 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  L0Memory_25 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  L0Memory_26 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  L0Memory_27 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  L0Memory_28 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  L0Memory_29 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  L0Memory_30 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  L0Memory_31 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  L0Memory_32 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  L0Memory_33 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  L0Memory_34 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  L0Memory_35 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  L0Memory_36 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  L0Memory_37 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  L0Memory_38 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  L0Memory_39 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  L0Memory_40 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  L0Memory_41 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  L0Memory_42 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  L0Memory_43 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  L0Memory_44 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  L0Memory_45 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  L0Memory_46 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  L0Memory_47 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  L0Memory_48 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  L0Memory_49 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  L0Memory_50 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  L0Memory_51 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  L0Memory_52 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  L0Memory_53 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  L0Memory_54 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  L0Memory_55 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  L0Memory_56 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  L0Memory_57 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  L0Memory_58 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  L0Memory_59 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  L0Memory_60 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  L0Memory_61 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  L0Memory_62 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  L0Memory_63 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  L0Memory_64 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  L0Memory_65 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  L0Memory_66 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  L0Memory_67 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  L0Memory_68 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  L0Memory_69 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  L0Memory_70 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  L0Memory_71 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  L0Memory_72 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  L0Memory_73 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  L0Memory_74 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  L0Memory_75 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  L0Memory_76 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  L0Memory_77 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  L0Memory_78 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  L0Memory_79 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  L0Memory_80 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  L0Memory_81 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  L0Memory_82 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  L0Memory_83 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  L0Memory_84 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  L0Memory_85 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  L0Memory_86 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  L0Memory_87 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  L0Memory_88 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  L0Memory_89 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  L0Memory_90 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  L0Memory_91 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  L0Memory_92 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  L0Memory_93 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  L0Memory_94 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  L0Memory_95 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  L0Memory_96 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  L0Memory_97 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  L0Memory_98 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  L0Memory_99 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  state = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  mux2out_reg = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  mux3out_reg = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  count = _RAND_104[9:0];
  _RAND_105 = {1{`RANDOM}};
  count_max = _RAND_105[9:0];
  _RAND_106 = {1{`RANDOM}};
  L0index_begin = _RAND_106[5:0];
  _RAND_107 = {1{`RANDOM}};
  GRU_out_width = _RAND_107[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PEArray(
  input         clock,
  input         reset,
  input  [15:0] io_From_above_0,
  input  [15:0] io_From_above_1,
  input  [15:0] io_From_above_2,
  input  [15:0] io_From_above_3,
  input  [15:0] io_From_above_4,
  input  [15:0] io_From_above_5,
  input  [15:0] io_From_above_6,
  input  [15:0] io_From_above_7,
  input  [15:0] io_From_above_8,
  input  [15:0] io_From_above_9,
  input  [15:0] io_From_above_10,
  input  [15:0] io_From_above_11,
  input  [11:0] io_PE_control_0_mask,
  input  [11:0] io_PE_control_1_mask,
  input  [2:0]  io_PE_control_2_control,
  input  [9:0]  io_PE_control_2_count,
  input  [5:0]  io_PE_control_2_L0index,
  input  [11:0] io_PE_control_2_mask,
  input  [7:0]  io_PE_control_2_gru_out_width,
  input  [3:0]  io_rd_data_mux,
  output [15:0] io_To_below_0,
  output [15:0] io_To_below_1,
  output [15:0] io_To_below_2,
  output [15:0] io_To_below_3,
  output [15:0] io_To_below_4,
  output [15:0] io_To_below_5,
  output [15:0] io_To_below_6,
  output [15:0] io_To_below_7,
  output [15:0] io_To_below_8,
  output [15:0] io_To_below_9,
  output [15:0] io_To_below_10,
  output [15:0] io_To_below_11,
  output [15:0] io_To_right_2
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  PE_Array_0_0_clock; // @[PEArray.scala 266:22]
  wire  PE_Array_0_0_reset; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_0_0_io_FromAbovePE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_0_0_io_FromL1; // @[PEArray.scala 266:22]
  wire [11:0] PE_Array_0_0_io_control_signal_mask; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_0_0_io_ToRightPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_0_0_io_ToBelowPE; // @[PEArray.scala 266:22]
  wire  PE_Array_0_1_clock; // @[PEArray.scala 266:22]
  wire  PE_Array_0_1_reset; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_0_1_io_FromAbovePE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_0_1_io_FromL1; // @[PEArray.scala 266:22]
  wire [11:0] PE_Array_0_1_io_control_signal_mask; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_0_1_io_ToRightPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_0_1_io_ToBelowPE; // @[PEArray.scala 266:22]
  wire  PE_Array_0_2_clock; // @[PEArray.scala 266:22]
  wire  PE_Array_0_2_reset; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_0_2_io_FromAbovePE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_0_2_io_FromL1; // @[PEArray.scala 266:22]
  wire [2:0] PE_Array_0_2_io_control_signal_control; // @[PEArray.scala 266:22]
  wire [9:0] PE_Array_0_2_io_control_signal_count; // @[PEArray.scala 266:22]
  wire [5:0] PE_Array_0_2_io_control_signal_L0index; // @[PEArray.scala 266:22]
  wire [11:0] PE_Array_0_2_io_control_signal_mask; // @[PEArray.scala 266:22]
  wire [7:0] PE_Array_0_2_io_control_signal_gru_out_width; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_0_2_io_ToRightPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_0_2_io_ToBelowPE; // @[PEArray.scala 266:22]
  wire  PE_Array_1_0_clock; // @[PEArray.scala 266:22]
  wire  PE_Array_1_0_reset; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_1_0_io_FromAbovePE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_1_0_io_FromLeftPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_1_0_io_FromL1; // @[PEArray.scala 266:22]
  wire [11:0] PE_Array_1_0_io_control_signal_mask; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_1_0_io_ToRightPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_1_0_io_ToBelowPE; // @[PEArray.scala 266:22]
  wire  PE_Array_1_1_clock; // @[PEArray.scala 266:22]
  wire  PE_Array_1_1_reset; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_1_1_io_FromAbovePE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_1_1_io_FromLeftPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_1_1_io_FromL1; // @[PEArray.scala 266:22]
  wire [11:0] PE_Array_1_1_io_control_signal_mask; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_1_1_io_ToRightPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_1_1_io_ToBelowPE; // @[PEArray.scala 266:22]
  wire  PE_Array_1_2_clock; // @[PEArray.scala 266:22]
  wire  PE_Array_1_2_reset; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_1_2_io_FromAbovePE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_1_2_io_FromLeftPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_1_2_io_FromL1; // @[PEArray.scala 266:22]
  wire [2:0] PE_Array_1_2_io_control_signal_control; // @[PEArray.scala 266:22]
  wire [9:0] PE_Array_1_2_io_control_signal_count; // @[PEArray.scala 266:22]
  wire [5:0] PE_Array_1_2_io_control_signal_L0index; // @[PEArray.scala 266:22]
  wire [11:0] PE_Array_1_2_io_control_signal_mask; // @[PEArray.scala 266:22]
  wire [7:0] PE_Array_1_2_io_control_signal_gru_out_width; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_1_2_io_ToRightPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_1_2_io_ToBelowPE; // @[PEArray.scala 266:22]
  wire  PE_Array_2_0_clock; // @[PEArray.scala 266:22]
  wire  PE_Array_2_0_reset; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_2_0_io_FromAbovePE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_2_0_io_FromLeftPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_2_0_io_FromL1; // @[PEArray.scala 266:22]
  wire [11:0] PE_Array_2_0_io_control_signal_mask; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_2_0_io_ToRightPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_2_0_io_ToBelowPE; // @[PEArray.scala 266:22]
  wire  PE_Array_2_1_clock; // @[PEArray.scala 266:22]
  wire  PE_Array_2_1_reset; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_2_1_io_FromAbovePE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_2_1_io_FromLeftPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_2_1_io_FromL1; // @[PEArray.scala 266:22]
  wire [11:0] PE_Array_2_1_io_control_signal_mask; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_2_1_io_ToRightPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_2_1_io_ToBelowPE; // @[PEArray.scala 266:22]
  wire  PE_Array_2_2_clock; // @[PEArray.scala 266:22]
  wire  PE_Array_2_2_reset; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_2_2_io_FromAbovePE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_2_2_io_FromLeftPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_2_2_io_FromL1; // @[PEArray.scala 266:22]
  wire [2:0] PE_Array_2_2_io_control_signal_control; // @[PEArray.scala 266:22]
  wire [9:0] PE_Array_2_2_io_control_signal_count; // @[PEArray.scala 266:22]
  wire [5:0] PE_Array_2_2_io_control_signal_L0index; // @[PEArray.scala 266:22]
  wire [11:0] PE_Array_2_2_io_control_signal_mask; // @[PEArray.scala 266:22]
  wire [7:0] PE_Array_2_2_io_control_signal_gru_out_width; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_2_2_io_ToRightPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_2_2_io_ToBelowPE; // @[PEArray.scala 266:22]
  wire  PE_Array_3_0_clock; // @[PEArray.scala 266:22]
  wire  PE_Array_3_0_reset; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_3_0_io_FromAbovePE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_3_0_io_FromLeftPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_3_0_io_FromL1; // @[PEArray.scala 266:22]
  wire [11:0] PE_Array_3_0_io_control_signal_mask; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_3_0_io_ToRightPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_3_0_io_ToBelowPE; // @[PEArray.scala 266:22]
  wire  PE_Array_3_1_clock; // @[PEArray.scala 266:22]
  wire  PE_Array_3_1_reset; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_3_1_io_FromAbovePE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_3_1_io_FromLeftPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_3_1_io_FromL1; // @[PEArray.scala 266:22]
  wire [11:0] PE_Array_3_1_io_control_signal_mask; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_3_1_io_ToRightPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_3_1_io_ToBelowPE; // @[PEArray.scala 266:22]
  wire  PE_Array_3_2_clock; // @[PEArray.scala 266:22]
  wire  PE_Array_3_2_reset; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_3_2_io_FromAbovePE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_3_2_io_FromLeftPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_3_2_io_FromL1; // @[PEArray.scala 266:22]
  wire [2:0] PE_Array_3_2_io_control_signal_control; // @[PEArray.scala 266:22]
  wire [9:0] PE_Array_3_2_io_control_signal_count; // @[PEArray.scala 266:22]
  wire [5:0] PE_Array_3_2_io_control_signal_L0index; // @[PEArray.scala 266:22]
  wire [11:0] PE_Array_3_2_io_control_signal_mask; // @[PEArray.scala 266:22]
  wire [7:0] PE_Array_3_2_io_control_signal_gru_out_width; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_3_2_io_ToRightPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_3_2_io_ToBelowPE; // @[PEArray.scala 266:22]
  wire  PE_Array_4_0_clock; // @[PEArray.scala 266:22]
  wire  PE_Array_4_0_reset; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_4_0_io_FromAbovePE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_4_0_io_FromLeftPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_4_0_io_FromL1; // @[PEArray.scala 266:22]
  wire [11:0] PE_Array_4_0_io_control_signal_mask; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_4_0_io_ToRightPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_4_0_io_ToBelowPE; // @[PEArray.scala 266:22]
  wire  PE_Array_4_1_clock; // @[PEArray.scala 266:22]
  wire  PE_Array_4_1_reset; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_4_1_io_FromAbovePE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_4_1_io_FromLeftPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_4_1_io_FromL1; // @[PEArray.scala 266:22]
  wire [11:0] PE_Array_4_1_io_control_signal_mask; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_4_1_io_ToRightPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_4_1_io_ToBelowPE; // @[PEArray.scala 266:22]
  wire  PE_Array_4_2_clock; // @[PEArray.scala 266:22]
  wire  PE_Array_4_2_reset; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_4_2_io_FromAbovePE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_4_2_io_FromLeftPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_4_2_io_FromL1; // @[PEArray.scala 266:22]
  wire [2:0] PE_Array_4_2_io_control_signal_control; // @[PEArray.scala 266:22]
  wire [9:0] PE_Array_4_2_io_control_signal_count; // @[PEArray.scala 266:22]
  wire [5:0] PE_Array_4_2_io_control_signal_L0index; // @[PEArray.scala 266:22]
  wire [11:0] PE_Array_4_2_io_control_signal_mask; // @[PEArray.scala 266:22]
  wire [7:0] PE_Array_4_2_io_control_signal_gru_out_width; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_4_2_io_ToRightPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_4_2_io_ToBelowPE; // @[PEArray.scala 266:22]
  wire  PE_Array_5_0_clock; // @[PEArray.scala 266:22]
  wire  PE_Array_5_0_reset; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_5_0_io_FromAbovePE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_5_0_io_FromLeftPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_5_0_io_FromL1; // @[PEArray.scala 266:22]
  wire [11:0] PE_Array_5_0_io_control_signal_mask; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_5_0_io_ToRightPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_5_0_io_ToBelowPE; // @[PEArray.scala 266:22]
  wire  PE_Array_5_1_clock; // @[PEArray.scala 266:22]
  wire  PE_Array_5_1_reset; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_5_1_io_FromAbovePE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_5_1_io_FromLeftPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_5_1_io_FromL1; // @[PEArray.scala 266:22]
  wire [11:0] PE_Array_5_1_io_control_signal_mask; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_5_1_io_ToRightPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_5_1_io_ToBelowPE; // @[PEArray.scala 266:22]
  wire  PE_Array_5_2_clock; // @[PEArray.scala 266:22]
  wire  PE_Array_5_2_reset; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_5_2_io_FromAbovePE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_5_2_io_FromLeftPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_5_2_io_FromL1; // @[PEArray.scala 266:22]
  wire [2:0] PE_Array_5_2_io_control_signal_control; // @[PEArray.scala 266:22]
  wire [9:0] PE_Array_5_2_io_control_signal_count; // @[PEArray.scala 266:22]
  wire [5:0] PE_Array_5_2_io_control_signal_L0index; // @[PEArray.scala 266:22]
  wire [11:0] PE_Array_5_2_io_control_signal_mask; // @[PEArray.scala 266:22]
  wire [7:0] PE_Array_5_2_io_control_signal_gru_out_width; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_5_2_io_ToRightPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_5_2_io_ToBelowPE; // @[PEArray.scala 266:22]
  wire  PE_Array_6_0_clock; // @[PEArray.scala 266:22]
  wire  PE_Array_6_0_reset; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_6_0_io_FromAbovePE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_6_0_io_FromLeftPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_6_0_io_FromL1; // @[PEArray.scala 266:22]
  wire [11:0] PE_Array_6_0_io_control_signal_mask; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_6_0_io_ToRightPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_6_0_io_ToBelowPE; // @[PEArray.scala 266:22]
  wire  PE_Array_6_1_clock; // @[PEArray.scala 266:22]
  wire  PE_Array_6_1_reset; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_6_1_io_FromAbovePE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_6_1_io_FromLeftPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_6_1_io_FromL1; // @[PEArray.scala 266:22]
  wire [11:0] PE_Array_6_1_io_control_signal_mask; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_6_1_io_ToRightPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_6_1_io_ToBelowPE; // @[PEArray.scala 266:22]
  wire  PE_Array_6_2_clock; // @[PEArray.scala 266:22]
  wire  PE_Array_6_2_reset; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_6_2_io_FromAbovePE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_6_2_io_FromLeftPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_6_2_io_FromL1; // @[PEArray.scala 266:22]
  wire [2:0] PE_Array_6_2_io_control_signal_control; // @[PEArray.scala 266:22]
  wire [9:0] PE_Array_6_2_io_control_signal_count; // @[PEArray.scala 266:22]
  wire [5:0] PE_Array_6_2_io_control_signal_L0index; // @[PEArray.scala 266:22]
  wire [11:0] PE_Array_6_2_io_control_signal_mask; // @[PEArray.scala 266:22]
  wire [7:0] PE_Array_6_2_io_control_signal_gru_out_width; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_6_2_io_ToRightPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_6_2_io_ToBelowPE; // @[PEArray.scala 266:22]
  wire  PE_Array_7_0_clock; // @[PEArray.scala 266:22]
  wire  PE_Array_7_0_reset; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_7_0_io_FromAbovePE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_7_0_io_FromLeftPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_7_0_io_FromL1; // @[PEArray.scala 266:22]
  wire [11:0] PE_Array_7_0_io_control_signal_mask; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_7_0_io_ToRightPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_7_0_io_ToBelowPE; // @[PEArray.scala 266:22]
  wire  PE_Array_7_1_clock; // @[PEArray.scala 266:22]
  wire  PE_Array_7_1_reset; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_7_1_io_FromAbovePE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_7_1_io_FromLeftPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_7_1_io_FromL1; // @[PEArray.scala 266:22]
  wire [11:0] PE_Array_7_1_io_control_signal_mask; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_7_1_io_ToRightPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_7_1_io_ToBelowPE; // @[PEArray.scala 266:22]
  wire  PE_Array_7_2_clock; // @[PEArray.scala 266:22]
  wire  PE_Array_7_2_reset; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_7_2_io_FromAbovePE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_7_2_io_FromLeftPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_7_2_io_FromL1; // @[PEArray.scala 266:22]
  wire [2:0] PE_Array_7_2_io_control_signal_control; // @[PEArray.scala 266:22]
  wire [9:0] PE_Array_7_2_io_control_signal_count; // @[PEArray.scala 266:22]
  wire [5:0] PE_Array_7_2_io_control_signal_L0index; // @[PEArray.scala 266:22]
  wire [11:0] PE_Array_7_2_io_control_signal_mask; // @[PEArray.scala 266:22]
  wire [7:0] PE_Array_7_2_io_control_signal_gru_out_width; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_7_2_io_ToRightPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_7_2_io_ToBelowPE; // @[PEArray.scala 266:22]
  wire  PE_Array_8_0_clock; // @[PEArray.scala 266:22]
  wire  PE_Array_8_0_reset; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_8_0_io_FromAbovePE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_8_0_io_FromLeftPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_8_0_io_FromL1; // @[PEArray.scala 266:22]
  wire [11:0] PE_Array_8_0_io_control_signal_mask; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_8_0_io_ToRightPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_8_0_io_ToBelowPE; // @[PEArray.scala 266:22]
  wire  PE_Array_8_1_clock; // @[PEArray.scala 266:22]
  wire  PE_Array_8_1_reset; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_8_1_io_FromAbovePE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_8_1_io_FromLeftPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_8_1_io_FromL1; // @[PEArray.scala 266:22]
  wire [11:0] PE_Array_8_1_io_control_signal_mask; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_8_1_io_ToRightPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_8_1_io_ToBelowPE; // @[PEArray.scala 266:22]
  wire  PE_Array_8_2_clock; // @[PEArray.scala 266:22]
  wire  PE_Array_8_2_reset; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_8_2_io_FromAbovePE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_8_2_io_FromLeftPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_8_2_io_FromL1; // @[PEArray.scala 266:22]
  wire [2:0] PE_Array_8_2_io_control_signal_control; // @[PEArray.scala 266:22]
  wire [9:0] PE_Array_8_2_io_control_signal_count; // @[PEArray.scala 266:22]
  wire [5:0] PE_Array_8_2_io_control_signal_L0index; // @[PEArray.scala 266:22]
  wire [11:0] PE_Array_8_2_io_control_signal_mask; // @[PEArray.scala 266:22]
  wire [7:0] PE_Array_8_2_io_control_signal_gru_out_width; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_8_2_io_ToRightPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_8_2_io_ToBelowPE; // @[PEArray.scala 266:22]
  wire  PE_Array_9_0_clock; // @[PEArray.scala 266:22]
  wire  PE_Array_9_0_reset; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_9_0_io_FromAbovePE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_9_0_io_FromLeftPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_9_0_io_FromL1; // @[PEArray.scala 266:22]
  wire [11:0] PE_Array_9_0_io_control_signal_mask; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_9_0_io_ToRightPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_9_0_io_ToBelowPE; // @[PEArray.scala 266:22]
  wire  PE_Array_9_1_clock; // @[PEArray.scala 266:22]
  wire  PE_Array_9_1_reset; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_9_1_io_FromAbovePE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_9_1_io_FromLeftPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_9_1_io_FromL1; // @[PEArray.scala 266:22]
  wire [11:0] PE_Array_9_1_io_control_signal_mask; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_9_1_io_ToRightPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_9_1_io_ToBelowPE; // @[PEArray.scala 266:22]
  wire  PE_Array_9_2_clock; // @[PEArray.scala 266:22]
  wire  PE_Array_9_2_reset; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_9_2_io_FromAbovePE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_9_2_io_FromLeftPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_9_2_io_FromL1; // @[PEArray.scala 266:22]
  wire [2:0] PE_Array_9_2_io_control_signal_control; // @[PEArray.scala 266:22]
  wire [9:0] PE_Array_9_2_io_control_signal_count; // @[PEArray.scala 266:22]
  wire [5:0] PE_Array_9_2_io_control_signal_L0index; // @[PEArray.scala 266:22]
  wire [11:0] PE_Array_9_2_io_control_signal_mask; // @[PEArray.scala 266:22]
  wire [7:0] PE_Array_9_2_io_control_signal_gru_out_width; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_9_2_io_ToRightPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_9_2_io_ToBelowPE; // @[PEArray.scala 266:22]
  wire  PE_Array_10_0_clock; // @[PEArray.scala 266:22]
  wire  PE_Array_10_0_reset; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_10_0_io_FromAbovePE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_10_0_io_FromLeftPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_10_0_io_FromL1; // @[PEArray.scala 266:22]
  wire [11:0] PE_Array_10_0_io_control_signal_mask; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_10_0_io_ToRightPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_10_0_io_ToBelowPE; // @[PEArray.scala 266:22]
  wire  PE_Array_10_1_clock; // @[PEArray.scala 266:22]
  wire  PE_Array_10_1_reset; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_10_1_io_FromAbovePE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_10_1_io_FromLeftPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_10_1_io_FromL1; // @[PEArray.scala 266:22]
  wire [11:0] PE_Array_10_1_io_control_signal_mask; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_10_1_io_ToRightPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_10_1_io_ToBelowPE; // @[PEArray.scala 266:22]
  wire  PE_Array_10_2_clock; // @[PEArray.scala 266:22]
  wire  PE_Array_10_2_reset; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_10_2_io_FromAbovePE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_10_2_io_FromLeftPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_10_2_io_FromL1; // @[PEArray.scala 266:22]
  wire [2:0] PE_Array_10_2_io_control_signal_control; // @[PEArray.scala 266:22]
  wire [9:0] PE_Array_10_2_io_control_signal_count; // @[PEArray.scala 266:22]
  wire [5:0] PE_Array_10_2_io_control_signal_L0index; // @[PEArray.scala 266:22]
  wire [11:0] PE_Array_10_2_io_control_signal_mask; // @[PEArray.scala 266:22]
  wire [7:0] PE_Array_10_2_io_control_signal_gru_out_width; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_10_2_io_ToRightPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_10_2_io_ToBelowPE; // @[PEArray.scala 266:22]
  wire  PE_Array_11_0_clock; // @[PEArray.scala 266:22]
  wire  PE_Array_11_0_reset; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_11_0_io_FromAbovePE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_11_0_io_FromLeftPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_11_0_io_FromL1; // @[PEArray.scala 266:22]
  wire [11:0] PE_Array_11_0_io_control_signal_mask; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_11_0_io_ToBelowPE; // @[PEArray.scala 266:22]
  wire  PE_Array_11_1_clock; // @[PEArray.scala 266:22]
  wire  PE_Array_11_1_reset; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_11_1_io_FromAbovePE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_11_1_io_FromLeftPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_11_1_io_FromL1; // @[PEArray.scala 266:22]
  wire [11:0] PE_Array_11_1_io_control_signal_mask; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_11_1_io_ToBelowPE; // @[PEArray.scala 266:22]
  wire  PE_Array_11_2_clock; // @[PEArray.scala 266:22]
  wire  PE_Array_11_2_reset; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_11_2_io_FromAbovePE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_11_2_io_FromLeftPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_11_2_io_FromL1; // @[PEArray.scala 266:22]
  wire [2:0] PE_Array_11_2_io_control_signal_control; // @[PEArray.scala 266:22]
  wire [9:0] PE_Array_11_2_io_control_signal_count; // @[PEArray.scala 266:22]
  wire [5:0] PE_Array_11_2_io_control_signal_L0index; // @[PEArray.scala 266:22]
  wire [11:0] PE_Array_11_2_io_control_signal_mask; // @[PEArray.scala 266:22]
  wire [7:0] PE_Array_11_2_io_control_signal_gru_out_width; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_11_2_io_ToRightPE; // @[PEArray.scala 266:22]
  wire [15:0] PE_Array_11_2_io_ToBelowPE; // @[PEArray.scala 266:22]
  reg [3:0] rd_data_mux_delay; // @[PEArray.scala 304:34]
  wire [15:0] _GEN_1 = 4'h1 == rd_data_mux_delay ? io_From_above_1 : io_From_above_0; // @[PEArray.scala 305:28 PEArray.scala 305:28]
  wire [15:0] _GEN_2 = 4'h2 == rd_data_mux_delay ? io_From_above_2 : _GEN_1; // @[PEArray.scala 305:28 PEArray.scala 305:28]
  wire [15:0] _GEN_3 = 4'h3 == rd_data_mux_delay ? io_From_above_3 : _GEN_2; // @[PEArray.scala 305:28 PEArray.scala 305:28]
  wire [15:0] _GEN_4 = 4'h4 == rd_data_mux_delay ? io_From_above_4 : _GEN_3; // @[PEArray.scala 305:28 PEArray.scala 305:28]
  wire [15:0] _GEN_5 = 4'h5 == rd_data_mux_delay ? io_From_above_5 : _GEN_4; // @[PEArray.scala 305:28 PEArray.scala 305:28]
  wire [15:0] _GEN_6 = 4'h6 == rd_data_mux_delay ? io_From_above_6 : _GEN_5; // @[PEArray.scala 305:28 PEArray.scala 305:28]
  wire [15:0] _GEN_7 = 4'h7 == rd_data_mux_delay ? io_From_above_7 : _GEN_6; // @[PEArray.scala 305:28 PEArray.scala 305:28]
  wire [15:0] _GEN_8 = 4'h8 == rd_data_mux_delay ? io_From_above_8 : _GEN_7; // @[PEArray.scala 305:28 PEArray.scala 305:28]
  wire [15:0] _GEN_9 = 4'h9 == rd_data_mux_delay ? io_From_above_9 : _GEN_8; // @[PEArray.scala 305:28 PEArray.scala 305:28]
  wire [15:0] _GEN_10 = 4'ha == rd_data_mux_delay ? io_From_above_10 : _GEN_9; // @[PEArray.scala 305:28 PEArray.scala 305:28]
  PE PE_Array_0_0 ( // @[PEArray.scala 266:22]
    .clock(PE_Array_0_0_clock),
    .reset(PE_Array_0_0_reset),
    .io_FromAbovePE(PE_Array_0_0_io_FromAbovePE),
    .io_FromL1(PE_Array_0_0_io_FromL1),
    .io_control_signal_mask(PE_Array_0_0_io_control_signal_mask),
    .io_ToRightPE(PE_Array_0_0_io_ToRightPE),
    .io_ToBelowPE(PE_Array_0_0_io_ToBelowPE)
  );
  PE_1 PE_Array_0_1 ( // @[PEArray.scala 266:22]
    .clock(PE_Array_0_1_clock),
    .reset(PE_Array_0_1_reset),
    .io_FromAbovePE(PE_Array_0_1_io_FromAbovePE),
    .io_FromL1(PE_Array_0_1_io_FromL1),
    .io_control_signal_mask(PE_Array_0_1_io_control_signal_mask),
    .io_ToRightPE(PE_Array_0_1_io_ToRightPE),
    .io_ToBelowPE(PE_Array_0_1_io_ToBelowPE)
  );
  PE_2 PE_Array_0_2 ( // @[PEArray.scala 266:22]
    .clock(PE_Array_0_2_clock),
    .reset(PE_Array_0_2_reset),
    .io_FromAbovePE(PE_Array_0_2_io_FromAbovePE),
    .io_FromL1(PE_Array_0_2_io_FromL1),
    .io_control_signal_control(PE_Array_0_2_io_control_signal_control),
    .io_control_signal_count(PE_Array_0_2_io_control_signal_count),
    .io_control_signal_L0index(PE_Array_0_2_io_control_signal_L0index),
    .io_control_signal_mask(PE_Array_0_2_io_control_signal_mask),
    .io_control_signal_gru_out_width(PE_Array_0_2_io_control_signal_gru_out_width),
    .io_ToRightPE(PE_Array_0_2_io_ToRightPE),
    .io_ToBelowPE(PE_Array_0_2_io_ToBelowPE)
  );
  PE_3 PE_Array_1_0 ( // @[PEArray.scala 266:22]
    .clock(PE_Array_1_0_clock),
    .reset(PE_Array_1_0_reset),
    .io_FromAbovePE(PE_Array_1_0_io_FromAbovePE),
    .io_FromLeftPE(PE_Array_1_0_io_FromLeftPE),
    .io_FromL1(PE_Array_1_0_io_FromL1),
    .io_control_signal_mask(PE_Array_1_0_io_control_signal_mask),
    .io_ToRightPE(PE_Array_1_0_io_ToRightPE),
    .io_ToBelowPE(PE_Array_1_0_io_ToBelowPE)
  );
  PE_4 PE_Array_1_1 ( // @[PEArray.scala 266:22]
    .clock(PE_Array_1_1_clock),
    .reset(PE_Array_1_1_reset),
    .io_FromAbovePE(PE_Array_1_1_io_FromAbovePE),
    .io_FromLeftPE(PE_Array_1_1_io_FromLeftPE),
    .io_FromL1(PE_Array_1_1_io_FromL1),
    .io_control_signal_mask(PE_Array_1_1_io_control_signal_mask),
    .io_ToRightPE(PE_Array_1_1_io_ToRightPE),
    .io_ToBelowPE(PE_Array_1_1_io_ToBelowPE)
  );
  PE_5 PE_Array_1_2 ( // @[PEArray.scala 266:22]
    .clock(PE_Array_1_2_clock),
    .reset(PE_Array_1_2_reset),
    .io_FromAbovePE(PE_Array_1_2_io_FromAbovePE),
    .io_FromLeftPE(PE_Array_1_2_io_FromLeftPE),
    .io_FromL1(PE_Array_1_2_io_FromL1),
    .io_control_signal_control(PE_Array_1_2_io_control_signal_control),
    .io_control_signal_count(PE_Array_1_2_io_control_signal_count),
    .io_control_signal_L0index(PE_Array_1_2_io_control_signal_L0index),
    .io_control_signal_mask(PE_Array_1_2_io_control_signal_mask),
    .io_control_signal_gru_out_width(PE_Array_1_2_io_control_signal_gru_out_width),
    .io_ToRightPE(PE_Array_1_2_io_ToRightPE),
    .io_ToBelowPE(PE_Array_1_2_io_ToBelowPE)
  );
  PE_6 PE_Array_2_0 ( // @[PEArray.scala 266:22]
    .clock(PE_Array_2_0_clock),
    .reset(PE_Array_2_0_reset),
    .io_FromAbovePE(PE_Array_2_0_io_FromAbovePE),
    .io_FromLeftPE(PE_Array_2_0_io_FromLeftPE),
    .io_FromL1(PE_Array_2_0_io_FromL1),
    .io_control_signal_mask(PE_Array_2_0_io_control_signal_mask),
    .io_ToRightPE(PE_Array_2_0_io_ToRightPE),
    .io_ToBelowPE(PE_Array_2_0_io_ToBelowPE)
  );
  PE_7 PE_Array_2_1 ( // @[PEArray.scala 266:22]
    .clock(PE_Array_2_1_clock),
    .reset(PE_Array_2_1_reset),
    .io_FromAbovePE(PE_Array_2_1_io_FromAbovePE),
    .io_FromLeftPE(PE_Array_2_1_io_FromLeftPE),
    .io_FromL1(PE_Array_2_1_io_FromL1),
    .io_control_signal_mask(PE_Array_2_1_io_control_signal_mask),
    .io_ToRightPE(PE_Array_2_1_io_ToRightPE),
    .io_ToBelowPE(PE_Array_2_1_io_ToBelowPE)
  );
  PE_8 PE_Array_2_2 ( // @[PEArray.scala 266:22]
    .clock(PE_Array_2_2_clock),
    .reset(PE_Array_2_2_reset),
    .io_FromAbovePE(PE_Array_2_2_io_FromAbovePE),
    .io_FromLeftPE(PE_Array_2_2_io_FromLeftPE),
    .io_FromL1(PE_Array_2_2_io_FromL1),
    .io_control_signal_control(PE_Array_2_2_io_control_signal_control),
    .io_control_signal_count(PE_Array_2_2_io_control_signal_count),
    .io_control_signal_L0index(PE_Array_2_2_io_control_signal_L0index),
    .io_control_signal_mask(PE_Array_2_2_io_control_signal_mask),
    .io_control_signal_gru_out_width(PE_Array_2_2_io_control_signal_gru_out_width),
    .io_ToRightPE(PE_Array_2_2_io_ToRightPE),
    .io_ToBelowPE(PE_Array_2_2_io_ToBelowPE)
  );
  PE_9 PE_Array_3_0 ( // @[PEArray.scala 266:22]
    .clock(PE_Array_3_0_clock),
    .reset(PE_Array_3_0_reset),
    .io_FromAbovePE(PE_Array_3_0_io_FromAbovePE),
    .io_FromLeftPE(PE_Array_3_0_io_FromLeftPE),
    .io_FromL1(PE_Array_3_0_io_FromL1),
    .io_control_signal_mask(PE_Array_3_0_io_control_signal_mask),
    .io_ToRightPE(PE_Array_3_0_io_ToRightPE),
    .io_ToBelowPE(PE_Array_3_0_io_ToBelowPE)
  );
  PE_10 PE_Array_3_1 ( // @[PEArray.scala 266:22]
    .clock(PE_Array_3_1_clock),
    .reset(PE_Array_3_1_reset),
    .io_FromAbovePE(PE_Array_3_1_io_FromAbovePE),
    .io_FromLeftPE(PE_Array_3_1_io_FromLeftPE),
    .io_FromL1(PE_Array_3_1_io_FromL1),
    .io_control_signal_mask(PE_Array_3_1_io_control_signal_mask),
    .io_ToRightPE(PE_Array_3_1_io_ToRightPE),
    .io_ToBelowPE(PE_Array_3_1_io_ToBelowPE)
  );
  PE_11 PE_Array_3_2 ( // @[PEArray.scala 266:22]
    .clock(PE_Array_3_2_clock),
    .reset(PE_Array_3_2_reset),
    .io_FromAbovePE(PE_Array_3_2_io_FromAbovePE),
    .io_FromLeftPE(PE_Array_3_2_io_FromLeftPE),
    .io_FromL1(PE_Array_3_2_io_FromL1),
    .io_control_signal_control(PE_Array_3_2_io_control_signal_control),
    .io_control_signal_count(PE_Array_3_2_io_control_signal_count),
    .io_control_signal_L0index(PE_Array_3_2_io_control_signal_L0index),
    .io_control_signal_mask(PE_Array_3_2_io_control_signal_mask),
    .io_control_signal_gru_out_width(PE_Array_3_2_io_control_signal_gru_out_width),
    .io_ToRightPE(PE_Array_3_2_io_ToRightPE),
    .io_ToBelowPE(PE_Array_3_2_io_ToBelowPE)
  );
  PE_12 PE_Array_4_0 ( // @[PEArray.scala 266:22]
    .clock(PE_Array_4_0_clock),
    .reset(PE_Array_4_0_reset),
    .io_FromAbovePE(PE_Array_4_0_io_FromAbovePE),
    .io_FromLeftPE(PE_Array_4_0_io_FromLeftPE),
    .io_FromL1(PE_Array_4_0_io_FromL1),
    .io_control_signal_mask(PE_Array_4_0_io_control_signal_mask),
    .io_ToRightPE(PE_Array_4_0_io_ToRightPE),
    .io_ToBelowPE(PE_Array_4_0_io_ToBelowPE)
  );
  PE_13 PE_Array_4_1 ( // @[PEArray.scala 266:22]
    .clock(PE_Array_4_1_clock),
    .reset(PE_Array_4_1_reset),
    .io_FromAbovePE(PE_Array_4_1_io_FromAbovePE),
    .io_FromLeftPE(PE_Array_4_1_io_FromLeftPE),
    .io_FromL1(PE_Array_4_1_io_FromL1),
    .io_control_signal_mask(PE_Array_4_1_io_control_signal_mask),
    .io_ToRightPE(PE_Array_4_1_io_ToRightPE),
    .io_ToBelowPE(PE_Array_4_1_io_ToBelowPE)
  );
  PE_14 PE_Array_4_2 ( // @[PEArray.scala 266:22]
    .clock(PE_Array_4_2_clock),
    .reset(PE_Array_4_2_reset),
    .io_FromAbovePE(PE_Array_4_2_io_FromAbovePE),
    .io_FromLeftPE(PE_Array_4_2_io_FromLeftPE),
    .io_FromL1(PE_Array_4_2_io_FromL1),
    .io_control_signal_control(PE_Array_4_2_io_control_signal_control),
    .io_control_signal_count(PE_Array_4_2_io_control_signal_count),
    .io_control_signal_L0index(PE_Array_4_2_io_control_signal_L0index),
    .io_control_signal_mask(PE_Array_4_2_io_control_signal_mask),
    .io_control_signal_gru_out_width(PE_Array_4_2_io_control_signal_gru_out_width),
    .io_ToRightPE(PE_Array_4_2_io_ToRightPE),
    .io_ToBelowPE(PE_Array_4_2_io_ToBelowPE)
  );
  PE_15 PE_Array_5_0 ( // @[PEArray.scala 266:22]
    .clock(PE_Array_5_0_clock),
    .reset(PE_Array_5_0_reset),
    .io_FromAbovePE(PE_Array_5_0_io_FromAbovePE),
    .io_FromLeftPE(PE_Array_5_0_io_FromLeftPE),
    .io_FromL1(PE_Array_5_0_io_FromL1),
    .io_control_signal_mask(PE_Array_5_0_io_control_signal_mask),
    .io_ToRightPE(PE_Array_5_0_io_ToRightPE),
    .io_ToBelowPE(PE_Array_5_0_io_ToBelowPE)
  );
  PE_16 PE_Array_5_1 ( // @[PEArray.scala 266:22]
    .clock(PE_Array_5_1_clock),
    .reset(PE_Array_5_1_reset),
    .io_FromAbovePE(PE_Array_5_1_io_FromAbovePE),
    .io_FromLeftPE(PE_Array_5_1_io_FromLeftPE),
    .io_FromL1(PE_Array_5_1_io_FromL1),
    .io_control_signal_mask(PE_Array_5_1_io_control_signal_mask),
    .io_ToRightPE(PE_Array_5_1_io_ToRightPE),
    .io_ToBelowPE(PE_Array_5_1_io_ToBelowPE)
  );
  PE_17 PE_Array_5_2 ( // @[PEArray.scala 266:22]
    .clock(PE_Array_5_2_clock),
    .reset(PE_Array_5_2_reset),
    .io_FromAbovePE(PE_Array_5_2_io_FromAbovePE),
    .io_FromLeftPE(PE_Array_5_2_io_FromLeftPE),
    .io_FromL1(PE_Array_5_2_io_FromL1),
    .io_control_signal_control(PE_Array_5_2_io_control_signal_control),
    .io_control_signal_count(PE_Array_5_2_io_control_signal_count),
    .io_control_signal_L0index(PE_Array_5_2_io_control_signal_L0index),
    .io_control_signal_mask(PE_Array_5_2_io_control_signal_mask),
    .io_control_signal_gru_out_width(PE_Array_5_2_io_control_signal_gru_out_width),
    .io_ToRightPE(PE_Array_5_2_io_ToRightPE),
    .io_ToBelowPE(PE_Array_5_2_io_ToBelowPE)
  );
  PE_18 PE_Array_6_0 ( // @[PEArray.scala 266:22]
    .clock(PE_Array_6_0_clock),
    .reset(PE_Array_6_0_reset),
    .io_FromAbovePE(PE_Array_6_0_io_FromAbovePE),
    .io_FromLeftPE(PE_Array_6_0_io_FromLeftPE),
    .io_FromL1(PE_Array_6_0_io_FromL1),
    .io_control_signal_mask(PE_Array_6_0_io_control_signal_mask),
    .io_ToRightPE(PE_Array_6_0_io_ToRightPE),
    .io_ToBelowPE(PE_Array_6_0_io_ToBelowPE)
  );
  PE_19 PE_Array_6_1 ( // @[PEArray.scala 266:22]
    .clock(PE_Array_6_1_clock),
    .reset(PE_Array_6_1_reset),
    .io_FromAbovePE(PE_Array_6_1_io_FromAbovePE),
    .io_FromLeftPE(PE_Array_6_1_io_FromLeftPE),
    .io_FromL1(PE_Array_6_1_io_FromL1),
    .io_control_signal_mask(PE_Array_6_1_io_control_signal_mask),
    .io_ToRightPE(PE_Array_6_1_io_ToRightPE),
    .io_ToBelowPE(PE_Array_6_1_io_ToBelowPE)
  );
  PE_20 PE_Array_6_2 ( // @[PEArray.scala 266:22]
    .clock(PE_Array_6_2_clock),
    .reset(PE_Array_6_2_reset),
    .io_FromAbovePE(PE_Array_6_2_io_FromAbovePE),
    .io_FromLeftPE(PE_Array_6_2_io_FromLeftPE),
    .io_FromL1(PE_Array_6_2_io_FromL1),
    .io_control_signal_control(PE_Array_6_2_io_control_signal_control),
    .io_control_signal_count(PE_Array_6_2_io_control_signal_count),
    .io_control_signal_L0index(PE_Array_6_2_io_control_signal_L0index),
    .io_control_signal_mask(PE_Array_6_2_io_control_signal_mask),
    .io_control_signal_gru_out_width(PE_Array_6_2_io_control_signal_gru_out_width),
    .io_ToRightPE(PE_Array_6_2_io_ToRightPE),
    .io_ToBelowPE(PE_Array_6_2_io_ToBelowPE)
  );
  PE_21 PE_Array_7_0 ( // @[PEArray.scala 266:22]
    .clock(PE_Array_7_0_clock),
    .reset(PE_Array_7_0_reset),
    .io_FromAbovePE(PE_Array_7_0_io_FromAbovePE),
    .io_FromLeftPE(PE_Array_7_0_io_FromLeftPE),
    .io_FromL1(PE_Array_7_0_io_FromL1),
    .io_control_signal_mask(PE_Array_7_0_io_control_signal_mask),
    .io_ToRightPE(PE_Array_7_0_io_ToRightPE),
    .io_ToBelowPE(PE_Array_7_0_io_ToBelowPE)
  );
  PE_22 PE_Array_7_1 ( // @[PEArray.scala 266:22]
    .clock(PE_Array_7_1_clock),
    .reset(PE_Array_7_1_reset),
    .io_FromAbovePE(PE_Array_7_1_io_FromAbovePE),
    .io_FromLeftPE(PE_Array_7_1_io_FromLeftPE),
    .io_FromL1(PE_Array_7_1_io_FromL1),
    .io_control_signal_mask(PE_Array_7_1_io_control_signal_mask),
    .io_ToRightPE(PE_Array_7_1_io_ToRightPE),
    .io_ToBelowPE(PE_Array_7_1_io_ToBelowPE)
  );
  PE_23 PE_Array_7_2 ( // @[PEArray.scala 266:22]
    .clock(PE_Array_7_2_clock),
    .reset(PE_Array_7_2_reset),
    .io_FromAbovePE(PE_Array_7_2_io_FromAbovePE),
    .io_FromLeftPE(PE_Array_7_2_io_FromLeftPE),
    .io_FromL1(PE_Array_7_2_io_FromL1),
    .io_control_signal_control(PE_Array_7_2_io_control_signal_control),
    .io_control_signal_count(PE_Array_7_2_io_control_signal_count),
    .io_control_signal_L0index(PE_Array_7_2_io_control_signal_L0index),
    .io_control_signal_mask(PE_Array_7_2_io_control_signal_mask),
    .io_control_signal_gru_out_width(PE_Array_7_2_io_control_signal_gru_out_width),
    .io_ToRightPE(PE_Array_7_2_io_ToRightPE),
    .io_ToBelowPE(PE_Array_7_2_io_ToBelowPE)
  );
  PE_24 PE_Array_8_0 ( // @[PEArray.scala 266:22]
    .clock(PE_Array_8_0_clock),
    .reset(PE_Array_8_0_reset),
    .io_FromAbovePE(PE_Array_8_0_io_FromAbovePE),
    .io_FromLeftPE(PE_Array_8_0_io_FromLeftPE),
    .io_FromL1(PE_Array_8_0_io_FromL1),
    .io_control_signal_mask(PE_Array_8_0_io_control_signal_mask),
    .io_ToRightPE(PE_Array_8_0_io_ToRightPE),
    .io_ToBelowPE(PE_Array_8_0_io_ToBelowPE)
  );
  PE_25 PE_Array_8_1 ( // @[PEArray.scala 266:22]
    .clock(PE_Array_8_1_clock),
    .reset(PE_Array_8_1_reset),
    .io_FromAbovePE(PE_Array_8_1_io_FromAbovePE),
    .io_FromLeftPE(PE_Array_8_1_io_FromLeftPE),
    .io_FromL1(PE_Array_8_1_io_FromL1),
    .io_control_signal_mask(PE_Array_8_1_io_control_signal_mask),
    .io_ToRightPE(PE_Array_8_1_io_ToRightPE),
    .io_ToBelowPE(PE_Array_8_1_io_ToBelowPE)
  );
  PE_26 PE_Array_8_2 ( // @[PEArray.scala 266:22]
    .clock(PE_Array_8_2_clock),
    .reset(PE_Array_8_2_reset),
    .io_FromAbovePE(PE_Array_8_2_io_FromAbovePE),
    .io_FromLeftPE(PE_Array_8_2_io_FromLeftPE),
    .io_FromL1(PE_Array_8_2_io_FromL1),
    .io_control_signal_control(PE_Array_8_2_io_control_signal_control),
    .io_control_signal_count(PE_Array_8_2_io_control_signal_count),
    .io_control_signal_L0index(PE_Array_8_2_io_control_signal_L0index),
    .io_control_signal_mask(PE_Array_8_2_io_control_signal_mask),
    .io_control_signal_gru_out_width(PE_Array_8_2_io_control_signal_gru_out_width),
    .io_ToRightPE(PE_Array_8_2_io_ToRightPE),
    .io_ToBelowPE(PE_Array_8_2_io_ToBelowPE)
  );
  PE_27 PE_Array_9_0 ( // @[PEArray.scala 266:22]
    .clock(PE_Array_9_0_clock),
    .reset(PE_Array_9_0_reset),
    .io_FromAbovePE(PE_Array_9_0_io_FromAbovePE),
    .io_FromLeftPE(PE_Array_9_0_io_FromLeftPE),
    .io_FromL1(PE_Array_9_0_io_FromL1),
    .io_control_signal_mask(PE_Array_9_0_io_control_signal_mask),
    .io_ToRightPE(PE_Array_9_0_io_ToRightPE),
    .io_ToBelowPE(PE_Array_9_0_io_ToBelowPE)
  );
  PE_28 PE_Array_9_1 ( // @[PEArray.scala 266:22]
    .clock(PE_Array_9_1_clock),
    .reset(PE_Array_9_1_reset),
    .io_FromAbovePE(PE_Array_9_1_io_FromAbovePE),
    .io_FromLeftPE(PE_Array_9_1_io_FromLeftPE),
    .io_FromL1(PE_Array_9_1_io_FromL1),
    .io_control_signal_mask(PE_Array_9_1_io_control_signal_mask),
    .io_ToRightPE(PE_Array_9_1_io_ToRightPE),
    .io_ToBelowPE(PE_Array_9_1_io_ToBelowPE)
  );
  PE_29 PE_Array_9_2 ( // @[PEArray.scala 266:22]
    .clock(PE_Array_9_2_clock),
    .reset(PE_Array_9_2_reset),
    .io_FromAbovePE(PE_Array_9_2_io_FromAbovePE),
    .io_FromLeftPE(PE_Array_9_2_io_FromLeftPE),
    .io_FromL1(PE_Array_9_2_io_FromL1),
    .io_control_signal_control(PE_Array_9_2_io_control_signal_control),
    .io_control_signal_count(PE_Array_9_2_io_control_signal_count),
    .io_control_signal_L0index(PE_Array_9_2_io_control_signal_L0index),
    .io_control_signal_mask(PE_Array_9_2_io_control_signal_mask),
    .io_control_signal_gru_out_width(PE_Array_9_2_io_control_signal_gru_out_width),
    .io_ToRightPE(PE_Array_9_2_io_ToRightPE),
    .io_ToBelowPE(PE_Array_9_2_io_ToBelowPE)
  );
  PE_30 PE_Array_10_0 ( // @[PEArray.scala 266:22]
    .clock(PE_Array_10_0_clock),
    .reset(PE_Array_10_0_reset),
    .io_FromAbovePE(PE_Array_10_0_io_FromAbovePE),
    .io_FromLeftPE(PE_Array_10_0_io_FromLeftPE),
    .io_FromL1(PE_Array_10_0_io_FromL1),
    .io_control_signal_mask(PE_Array_10_0_io_control_signal_mask),
    .io_ToRightPE(PE_Array_10_0_io_ToRightPE),
    .io_ToBelowPE(PE_Array_10_0_io_ToBelowPE)
  );
  PE_31 PE_Array_10_1 ( // @[PEArray.scala 266:22]
    .clock(PE_Array_10_1_clock),
    .reset(PE_Array_10_1_reset),
    .io_FromAbovePE(PE_Array_10_1_io_FromAbovePE),
    .io_FromLeftPE(PE_Array_10_1_io_FromLeftPE),
    .io_FromL1(PE_Array_10_1_io_FromL1),
    .io_control_signal_mask(PE_Array_10_1_io_control_signal_mask),
    .io_ToRightPE(PE_Array_10_1_io_ToRightPE),
    .io_ToBelowPE(PE_Array_10_1_io_ToBelowPE)
  );
  PE_32 PE_Array_10_2 ( // @[PEArray.scala 266:22]
    .clock(PE_Array_10_2_clock),
    .reset(PE_Array_10_2_reset),
    .io_FromAbovePE(PE_Array_10_2_io_FromAbovePE),
    .io_FromLeftPE(PE_Array_10_2_io_FromLeftPE),
    .io_FromL1(PE_Array_10_2_io_FromL1),
    .io_control_signal_control(PE_Array_10_2_io_control_signal_control),
    .io_control_signal_count(PE_Array_10_2_io_control_signal_count),
    .io_control_signal_L0index(PE_Array_10_2_io_control_signal_L0index),
    .io_control_signal_mask(PE_Array_10_2_io_control_signal_mask),
    .io_control_signal_gru_out_width(PE_Array_10_2_io_control_signal_gru_out_width),
    .io_ToRightPE(PE_Array_10_2_io_ToRightPE),
    .io_ToBelowPE(PE_Array_10_2_io_ToBelowPE)
  );
  PE_33 PE_Array_11_0 ( // @[PEArray.scala 266:22]
    .clock(PE_Array_11_0_clock),
    .reset(PE_Array_11_0_reset),
    .io_FromAbovePE(PE_Array_11_0_io_FromAbovePE),
    .io_FromLeftPE(PE_Array_11_0_io_FromLeftPE),
    .io_FromL1(PE_Array_11_0_io_FromL1),
    .io_control_signal_mask(PE_Array_11_0_io_control_signal_mask),
    .io_ToBelowPE(PE_Array_11_0_io_ToBelowPE)
  );
  PE_34 PE_Array_11_1 ( // @[PEArray.scala 266:22]
    .clock(PE_Array_11_1_clock),
    .reset(PE_Array_11_1_reset),
    .io_FromAbovePE(PE_Array_11_1_io_FromAbovePE),
    .io_FromLeftPE(PE_Array_11_1_io_FromLeftPE),
    .io_FromL1(PE_Array_11_1_io_FromL1),
    .io_control_signal_mask(PE_Array_11_1_io_control_signal_mask),
    .io_ToBelowPE(PE_Array_11_1_io_ToBelowPE)
  );
  PE_35 PE_Array_11_2 ( // @[PEArray.scala 266:22]
    .clock(PE_Array_11_2_clock),
    .reset(PE_Array_11_2_reset),
    .io_FromAbovePE(PE_Array_11_2_io_FromAbovePE),
    .io_FromLeftPE(PE_Array_11_2_io_FromLeftPE),
    .io_FromL1(PE_Array_11_2_io_FromL1),
    .io_control_signal_control(PE_Array_11_2_io_control_signal_control),
    .io_control_signal_count(PE_Array_11_2_io_control_signal_count),
    .io_control_signal_L0index(PE_Array_11_2_io_control_signal_L0index),
    .io_control_signal_mask(PE_Array_11_2_io_control_signal_mask),
    .io_control_signal_gru_out_width(PE_Array_11_2_io_control_signal_gru_out_width),
    .io_ToRightPE(PE_Array_11_2_io_ToRightPE),
    .io_ToBelowPE(PE_Array_11_2_io_ToBelowPE)
  );
  assign io_To_below_0 = PE_Array_0_2_io_ToBelowPE; // @[PEArray.scala 298:20]
  assign io_To_below_1 = PE_Array_1_2_io_ToBelowPE; // @[PEArray.scala 298:20]
  assign io_To_below_2 = PE_Array_2_2_io_ToBelowPE; // @[PEArray.scala 298:20]
  assign io_To_below_3 = PE_Array_3_2_io_ToBelowPE; // @[PEArray.scala 298:20]
  assign io_To_below_4 = PE_Array_4_2_io_ToBelowPE; // @[PEArray.scala 298:20]
  assign io_To_below_5 = PE_Array_5_2_io_ToBelowPE; // @[PEArray.scala 298:20]
  assign io_To_below_6 = PE_Array_6_2_io_ToBelowPE; // @[PEArray.scala 298:20]
  assign io_To_below_7 = PE_Array_7_2_io_ToBelowPE; // @[PEArray.scala 298:20]
  assign io_To_below_8 = PE_Array_8_2_io_ToBelowPE; // @[PEArray.scala 298:20]
  assign io_To_below_9 = PE_Array_9_2_io_ToBelowPE; // @[PEArray.scala 298:20]
  assign io_To_below_10 = PE_Array_10_2_io_ToBelowPE; // @[PEArray.scala 298:20]
  assign io_To_below_11 = PE_Array_11_2_io_ToBelowPE; // @[PEArray.scala 298:20]
  assign io_To_right_2 = PE_Array_11_2_io_ToRightPE; // @[PEArray.scala 314:20]
  assign PE_Array_0_0_clock = clock;
  assign PE_Array_0_0_reset = reset;
  assign PE_Array_0_0_io_FromAbovePE = PE_Array_0_2_io_ToBelowPE; // @[PEArray.scala 297:35]
  assign PE_Array_0_0_io_FromL1 = io_From_above_0; // @[PEArray.scala 302:28]
  assign PE_Array_0_0_io_control_signal_mask = io_PE_control_0_mask; // @[PEArray.scala 274:40]
  assign PE_Array_0_1_clock = clock;
  assign PE_Array_0_1_reset = reset;
  assign PE_Array_0_1_io_FromAbovePE = PE_Array_0_0_io_ToBelowPE; // @[PEArray.scala 291:39]
  assign PE_Array_0_1_io_FromL1 = io_From_above_0; // @[PEArray.scala 303:28]
  assign PE_Array_0_1_io_control_signal_mask = io_PE_control_1_mask; // @[PEArray.scala 274:40]
  assign PE_Array_0_2_clock = clock;
  assign PE_Array_0_2_reset = reset;
  assign PE_Array_0_2_io_FromAbovePE = PE_Array_0_1_io_ToBelowPE; // @[PEArray.scala 291:39]
  assign PE_Array_0_2_io_FromL1 = 4'hb == rd_data_mux_delay ? io_From_above_11 : _GEN_10; // @[PEArray.scala 305:28 PEArray.scala 305:28]
  assign PE_Array_0_2_io_control_signal_control = io_PE_control_2_control; // @[PEArray.scala 274:40]
  assign PE_Array_0_2_io_control_signal_count = io_PE_control_2_count; // @[PEArray.scala 274:40]
  assign PE_Array_0_2_io_control_signal_L0index = io_PE_control_2_L0index; // @[PEArray.scala 274:40]
  assign PE_Array_0_2_io_control_signal_mask = io_PE_control_2_mask; // @[PEArray.scala 274:40]
  assign PE_Array_0_2_io_control_signal_gru_out_width = io_PE_control_2_gru_out_width; // @[PEArray.scala 274:40]
  assign PE_Array_1_0_clock = clock;
  assign PE_Array_1_0_reset = reset;
  assign PE_Array_1_0_io_FromAbovePE = PE_Array_1_2_io_ToBelowPE; // @[PEArray.scala 297:35]
  assign PE_Array_1_0_io_FromLeftPE = PE_Array_0_0_io_ToRightPE; // @[PEArray.scala 281:38]
  assign PE_Array_1_0_io_FromL1 = io_From_above_1; // @[PEArray.scala 308:32]
  assign PE_Array_1_0_io_control_signal_mask = io_PE_control_0_mask; // @[PEArray.scala 274:40]
  assign PE_Array_1_1_clock = clock;
  assign PE_Array_1_1_reset = reset;
  assign PE_Array_1_1_io_FromAbovePE = PE_Array_1_0_io_ToBelowPE; // @[PEArray.scala 291:39]
  assign PE_Array_1_1_io_FromLeftPE = PE_Array_0_1_io_ToRightPE; // @[PEArray.scala 281:38]
  assign PE_Array_1_1_io_FromL1 = io_From_above_1; // @[PEArray.scala 308:32]
  assign PE_Array_1_1_io_control_signal_mask = io_PE_control_1_mask; // @[PEArray.scala 274:40]
  assign PE_Array_1_2_clock = clock;
  assign PE_Array_1_2_reset = reset;
  assign PE_Array_1_2_io_FromAbovePE = PE_Array_1_1_io_ToBelowPE; // @[PEArray.scala 291:39]
  assign PE_Array_1_2_io_FromLeftPE = PE_Array_0_2_io_ToRightPE; // @[PEArray.scala 281:38]
  assign PE_Array_1_2_io_FromL1 = io_From_above_1; // @[PEArray.scala 308:32]
  assign PE_Array_1_2_io_control_signal_control = io_PE_control_2_control; // @[PEArray.scala 274:40]
  assign PE_Array_1_2_io_control_signal_count = io_PE_control_2_count; // @[PEArray.scala 274:40]
  assign PE_Array_1_2_io_control_signal_L0index = io_PE_control_2_L0index; // @[PEArray.scala 274:40]
  assign PE_Array_1_2_io_control_signal_mask = io_PE_control_2_mask; // @[PEArray.scala 274:40]
  assign PE_Array_1_2_io_control_signal_gru_out_width = io_PE_control_2_gru_out_width; // @[PEArray.scala 274:40]
  assign PE_Array_2_0_clock = clock;
  assign PE_Array_2_0_reset = reset;
  assign PE_Array_2_0_io_FromAbovePE = PE_Array_2_2_io_ToBelowPE; // @[PEArray.scala 297:35]
  assign PE_Array_2_0_io_FromLeftPE = PE_Array_1_0_io_ToRightPE; // @[PEArray.scala 281:38]
  assign PE_Array_2_0_io_FromL1 = io_From_above_2; // @[PEArray.scala 308:32]
  assign PE_Array_2_0_io_control_signal_mask = io_PE_control_0_mask; // @[PEArray.scala 274:40]
  assign PE_Array_2_1_clock = clock;
  assign PE_Array_2_1_reset = reset;
  assign PE_Array_2_1_io_FromAbovePE = PE_Array_2_0_io_ToBelowPE; // @[PEArray.scala 291:39]
  assign PE_Array_2_1_io_FromLeftPE = PE_Array_1_1_io_ToRightPE; // @[PEArray.scala 281:38]
  assign PE_Array_2_1_io_FromL1 = io_From_above_2; // @[PEArray.scala 308:32]
  assign PE_Array_2_1_io_control_signal_mask = io_PE_control_1_mask; // @[PEArray.scala 274:40]
  assign PE_Array_2_2_clock = clock;
  assign PE_Array_2_2_reset = reset;
  assign PE_Array_2_2_io_FromAbovePE = PE_Array_2_1_io_ToBelowPE; // @[PEArray.scala 291:39]
  assign PE_Array_2_2_io_FromLeftPE = PE_Array_1_2_io_ToRightPE; // @[PEArray.scala 281:38]
  assign PE_Array_2_2_io_FromL1 = io_From_above_2; // @[PEArray.scala 308:32]
  assign PE_Array_2_2_io_control_signal_control = io_PE_control_2_control; // @[PEArray.scala 274:40]
  assign PE_Array_2_2_io_control_signal_count = io_PE_control_2_count; // @[PEArray.scala 274:40]
  assign PE_Array_2_2_io_control_signal_L0index = io_PE_control_2_L0index; // @[PEArray.scala 274:40]
  assign PE_Array_2_2_io_control_signal_mask = io_PE_control_2_mask; // @[PEArray.scala 274:40]
  assign PE_Array_2_2_io_control_signal_gru_out_width = io_PE_control_2_gru_out_width; // @[PEArray.scala 274:40]
  assign PE_Array_3_0_clock = clock;
  assign PE_Array_3_0_reset = reset;
  assign PE_Array_3_0_io_FromAbovePE = PE_Array_3_2_io_ToBelowPE; // @[PEArray.scala 297:35]
  assign PE_Array_3_0_io_FromLeftPE = PE_Array_2_0_io_ToRightPE; // @[PEArray.scala 281:38]
  assign PE_Array_3_0_io_FromL1 = io_From_above_3; // @[PEArray.scala 308:32]
  assign PE_Array_3_0_io_control_signal_mask = io_PE_control_0_mask; // @[PEArray.scala 274:40]
  assign PE_Array_3_1_clock = clock;
  assign PE_Array_3_1_reset = reset;
  assign PE_Array_3_1_io_FromAbovePE = PE_Array_3_0_io_ToBelowPE; // @[PEArray.scala 291:39]
  assign PE_Array_3_1_io_FromLeftPE = PE_Array_2_1_io_ToRightPE; // @[PEArray.scala 281:38]
  assign PE_Array_3_1_io_FromL1 = io_From_above_3; // @[PEArray.scala 308:32]
  assign PE_Array_3_1_io_control_signal_mask = io_PE_control_1_mask; // @[PEArray.scala 274:40]
  assign PE_Array_3_2_clock = clock;
  assign PE_Array_3_2_reset = reset;
  assign PE_Array_3_2_io_FromAbovePE = PE_Array_3_1_io_ToBelowPE; // @[PEArray.scala 291:39]
  assign PE_Array_3_2_io_FromLeftPE = PE_Array_2_2_io_ToRightPE; // @[PEArray.scala 281:38]
  assign PE_Array_3_2_io_FromL1 = io_From_above_3; // @[PEArray.scala 308:32]
  assign PE_Array_3_2_io_control_signal_control = io_PE_control_2_control; // @[PEArray.scala 274:40]
  assign PE_Array_3_2_io_control_signal_count = io_PE_control_2_count; // @[PEArray.scala 274:40]
  assign PE_Array_3_2_io_control_signal_L0index = io_PE_control_2_L0index; // @[PEArray.scala 274:40]
  assign PE_Array_3_2_io_control_signal_mask = io_PE_control_2_mask; // @[PEArray.scala 274:40]
  assign PE_Array_3_2_io_control_signal_gru_out_width = io_PE_control_2_gru_out_width; // @[PEArray.scala 274:40]
  assign PE_Array_4_0_clock = clock;
  assign PE_Array_4_0_reset = reset;
  assign PE_Array_4_0_io_FromAbovePE = PE_Array_4_2_io_ToBelowPE; // @[PEArray.scala 297:35]
  assign PE_Array_4_0_io_FromLeftPE = PE_Array_3_0_io_ToRightPE; // @[PEArray.scala 281:38]
  assign PE_Array_4_0_io_FromL1 = io_From_above_4; // @[PEArray.scala 308:32]
  assign PE_Array_4_0_io_control_signal_mask = io_PE_control_0_mask; // @[PEArray.scala 274:40]
  assign PE_Array_4_1_clock = clock;
  assign PE_Array_4_1_reset = reset;
  assign PE_Array_4_1_io_FromAbovePE = PE_Array_4_0_io_ToBelowPE; // @[PEArray.scala 291:39]
  assign PE_Array_4_1_io_FromLeftPE = PE_Array_3_1_io_ToRightPE; // @[PEArray.scala 281:38]
  assign PE_Array_4_1_io_FromL1 = io_From_above_4; // @[PEArray.scala 308:32]
  assign PE_Array_4_1_io_control_signal_mask = io_PE_control_1_mask; // @[PEArray.scala 274:40]
  assign PE_Array_4_2_clock = clock;
  assign PE_Array_4_2_reset = reset;
  assign PE_Array_4_2_io_FromAbovePE = PE_Array_4_1_io_ToBelowPE; // @[PEArray.scala 291:39]
  assign PE_Array_4_2_io_FromLeftPE = PE_Array_3_2_io_ToRightPE; // @[PEArray.scala 281:38]
  assign PE_Array_4_2_io_FromL1 = io_From_above_4; // @[PEArray.scala 308:32]
  assign PE_Array_4_2_io_control_signal_control = io_PE_control_2_control; // @[PEArray.scala 274:40]
  assign PE_Array_4_2_io_control_signal_count = io_PE_control_2_count; // @[PEArray.scala 274:40]
  assign PE_Array_4_2_io_control_signal_L0index = io_PE_control_2_L0index; // @[PEArray.scala 274:40]
  assign PE_Array_4_2_io_control_signal_mask = io_PE_control_2_mask; // @[PEArray.scala 274:40]
  assign PE_Array_4_2_io_control_signal_gru_out_width = io_PE_control_2_gru_out_width; // @[PEArray.scala 274:40]
  assign PE_Array_5_0_clock = clock;
  assign PE_Array_5_0_reset = reset;
  assign PE_Array_5_0_io_FromAbovePE = PE_Array_5_2_io_ToBelowPE; // @[PEArray.scala 297:35]
  assign PE_Array_5_0_io_FromLeftPE = PE_Array_4_0_io_ToRightPE; // @[PEArray.scala 281:38]
  assign PE_Array_5_0_io_FromL1 = io_From_above_5; // @[PEArray.scala 308:32]
  assign PE_Array_5_0_io_control_signal_mask = io_PE_control_0_mask; // @[PEArray.scala 274:40]
  assign PE_Array_5_1_clock = clock;
  assign PE_Array_5_1_reset = reset;
  assign PE_Array_5_1_io_FromAbovePE = PE_Array_5_0_io_ToBelowPE; // @[PEArray.scala 291:39]
  assign PE_Array_5_1_io_FromLeftPE = PE_Array_4_1_io_ToRightPE; // @[PEArray.scala 281:38]
  assign PE_Array_5_1_io_FromL1 = io_From_above_5; // @[PEArray.scala 308:32]
  assign PE_Array_5_1_io_control_signal_mask = io_PE_control_1_mask; // @[PEArray.scala 274:40]
  assign PE_Array_5_2_clock = clock;
  assign PE_Array_5_2_reset = reset;
  assign PE_Array_5_2_io_FromAbovePE = PE_Array_5_1_io_ToBelowPE; // @[PEArray.scala 291:39]
  assign PE_Array_5_2_io_FromLeftPE = PE_Array_4_2_io_ToRightPE; // @[PEArray.scala 281:38]
  assign PE_Array_5_2_io_FromL1 = io_From_above_5; // @[PEArray.scala 308:32]
  assign PE_Array_5_2_io_control_signal_control = io_PE_control_2_control; // @[PEArray.scala 274:40]
  assign PE_Array_5_2_io_control_signal_count = io_PE_control_2_count; // @[PEArray.scala 274:40]
  assign PE_Array_5_2_io_control_signal_L0index = io_PE_control_2_L0index; // @[PEArray.scala 274:40]
  assign PE_Array_5_2_io_control_signal_mask = io_PE_control_2_mask; // @[PEArray.scala 274:40]
  assign PE_Array_5_2_io_control_signal_gru_out_width = io_PE_control_2_gru_out_width; // @[PEArray.scala 274:40]
  assign PE_Array_6_0_clock = clock;
  assign PE_Array_6_0_reset = reset;
  assign PE_Array_6_0_io_FromAbovePE = PE_Array_6_2_io_ToBelowPE; // @[PEArray.scala 297:35]
  assign PE_Array_6_0_io_FromLeftPE = PE_Array_5_0_io_ToRightPE; // @[PEArray.scala 281:38]
  assign PE_Array_6_0_io_FromL1 = io_From_above_6; // @[PEArray.scala 308:32]
  assign PE_Array_6_0_io_control_signal_mask = io_PE_control_0_mask; // @[PEArray.scala 274:40]
  assign PE_Array_6_1_clock = clock;
  assign PE_Array_6_1_reset = reset;
  assign PE_Array_6_1_io_FromAbovePE = PE_Array_6_0_io_ToBelowPE; // @[PEArray.scala 291:39]
  assign PE_Array_6_1_io_FromLeftPE = PE_Array_5_1_io_ToRightPE; // @[PEArray.scala 281:38]
  assign PE_Array_6_1_io_FromL1 = io_From_above_6; // @[PEArray.scala 308:32]
  assign PE_Array_6_1_io_control_signal_mask = io_PE_control_1_mask; // @[PEArray.scala 274:40]
  assign PE_Array_6_2_clock = clock;
  assign PE_Array_6_2_reset = reset;
  assign PE_Array_6_2_io_FromAbovePE = PE_Array_6_1_io_ToBelowPE; // @[PEArray.scala 291:39]
  assign PE_Array_6_2_io_FromLeftPE = PE_Array_5_2_io_ToRightPE; // @[PEArray.scala 281:38]
  assign PE_Array_6_2_io_FromL1 = io_From_above_6; // @[PEArray.scala 308:32]
  assign PE_Array_6_2_io_control_signal_control = io_PE_control_2_control; // @[PEArray.scala 274:40]
  assign PE_Array_6_2_io_control_signal_count = io_PE_control_2_count; // @[PEArray.scala 274:40]
  assign PE_Array_6_2_io_control_signal_L0index = io_PE_control_2_L0index; // @[PEArray.scala 274:40]
  assign PE_Array_6_2_io_control_signal_mask = io_PE_control_2_mask; // @[PEArray.scala 274:40]
  assign PE_Array_6_2_io_control_signal_gru_out_width = io_PE_control_2_gru_out_width; // @[PEArray.scala 274:40]
  assign PE_Array_7_0_clock = clock;
  assign PE_Array_7_0_reset = reset;
  assign PE_Array_7_0_io_FromAbovePE = PE_Array_7_2_io_ToBelowPE; // @[PEArray.scala 297:35]
  assign PE_Array_7_0_io_FromLeftPE = PE_Array_6_0_io_ToRightPE; // @[PEArray.scala 281:38]
  assign PE_Array_7_0_io_FromL1 = io_From_above_7; // @[PEArray.scala 308:32]
  assign PE_Array_7_0_io_control_signal_mask = io_PE_control_0_mask; // @[PEArray.scala 274:40]
  assign PE_Array_7_1_clock = clock;
  assign PE_Array_7_1_reset = reset;
  assign PE_Array_7_1_io_FromAbovePE = PE_Array_7_0_io_ToBelowPE; // @[PEArray.scala 291:39]
  assign PE_Array_7_1_io_FromLeftPE = PE_Array_6_1_io_ToRightPE; // @[PEArray.scala 281:38]
  assign PE_Array_7_1_io_FromL1 = io_From_above_7; // @[PEArray.scala 308:32]
  assign PE_Array_7_1_io_control_signal_mask = io_PE_control_1_mask; // @[PEArray.scala 274:40]
  assign PE_Array_7_2_clock = clock;
  assign PE_Array_7_2_reset = reset;
  assign PE_Array_7_2_io_FromAbovePE = PE_Array_7_1_io_ToBelowPE; // @[PEArray.scala 291:39]
  assign PE_Array_7_2_io_FromLeftPE = PE_Array_6_2_io_ToRightPE; // @[PEArray.scala 281:38]
  assign PE_Array_7_2_io_FromL1 = io_From_above_7; // @[PEArray.scala 308:32]
  assign PE_Array_7_2_io_control_signal_control = io_PE_control_2_control; // @[PEArray.scala 274:40]
  assign PE_Array_7_2_io_control_signal_count = io_PE_control_2_count; // @[PEArray.scala 274:40]
  assign PE_Array_7_2_io_control_signal_L0index = io_PE_control_2_L0index; // @[PEArray.scala 274:40]
  assign PE_Array_7_2_io_control_signal_mask = io_PE_control_2_mask; // @[PEArray.scala 274:40]
  assign PE_Array_7_2_io_control_signal_gru_out_width = io_PE_control_2_gru_out_width; // @[PEArray.scala 274:40]
  assign PE_Array_8_0_clock = clock;
  assign PE_Array_8_0_reset = reset;
  assign PE_Array_8_0_io_FromAbovePE = PE_Array_8_2_io_ToBelowPE; // @[PEArray.scala 297:35]
  assign PE_Array_8_0_io_FromLeftPE = PE_Array_7_0_io_ToRightPE; // @[PEArray.scala 281:38]
  assign PE_Array_8_0_io_FromL1 = io_From_above_8; // @[PEArray.scala 308:32]
  assign PE_Array_8_0_io_control_signal_mask = io_PE_control_0_mask; // @[PEArray.scala 274:40]
  assign PE_Array_8_1_clock = clock;
  assign PE_Array_8_1_reset = reset;
  assign PE_Array_8_1_io_FromAbovePE = PE_Array_8_0_io_ToBelowPE; // @[PEArray.scala 291:39]
  assign PE_Array_8_1_io_FromLeftPE = PE_Array_7_1_io_ToRightPE; // @[PEArray.scala 281:38]
  assign PE_Array_8_1_io_FromL1 = io_From_above_8; // @[PEArray.scala 308:32]
  assign PE_Array_8_1_io_control_signal_mask = io_PE_control_1_mask; // @[PEArray.scala 274:40]
  assign PE_Array_8_2_clock = clock;
  assign PE_Array_8_2_reset = reset;
  assign PE_Array_8_2_io_FromAbovePE = PE_Array_8_1_io_ToBelowPE; // @[PEArray.scala 291:39]
  assign PE_Array_8_2_io_FromLeftPE = PE_Array_7_2_io_ToRightPE; // @[PEArray.scala 281:38]
  assign PE_Array_8_2_io_FromL1 = io_From_above_8; // @[PEArray.scala 308:32]
  assign PE_Array_8_2_io_control_signal_control = io_PE_control_2_control; // @[PEArray.scala 274:40]
  assign PE_Array_8_2_io_control_signal_count = io_PE_control_2_count; // @[PEArray.scala 274:40]
  assign PE_Array_8_2_io_control_signal_L0index = io_PE_control_2_L0index; // @[PEArray.scala 274:40]
  assign PE_Array_8_2_io_control_signal_mask = io_PE_control_2_mask; // @[PEArray.scala 274:40]
  assign PE_Array_8_2_io_control_signal_gru_out_width = io_PE_control_2_gru_out_width; // @[PEArray.scala 274:40]
  assign PE_Array_9_0_clock = clock;
  assign PE_Array_9_0_reset = reset;
  assign PE_Array_9_0_io_FromAbovePE = PE_Array_9_2_io_ToBelowPE; // @[PEArray.scala 297:35]
  assign PE_Array_9_0_io_FromLeftPE = PE_Array_8_0_io_ToRightPE; // @[PEArray.scala 281:38]
  assign PE_Array_9_0_io_FromL1 = io_From_above_9; // @[PEArray.scala 308:32]
  assign PE_Array_9_0_io_control_signal_mask = io_PE_control_0_mask; // @[PEArray.scala 274:40]
  assign PE_Array_9_1_clock = clock;
  assign PE_Array_9_1_reset = reset;
  assign PE_Array_9_1_io_FromAbovePE = PE_Array_9_0_io_ToBelowPE; // @[PEArray.scala 291:39]
  assign PE_Array_9_1_io_FromLeftPE = PE_Array_8_1_io_ToRightPE; // @[PEArray.scala 281:38]
  assign PE_Array_9_1_io_FromL1 = io_From_above_9; // @[PEArray.scala 308:32]
  assign PE_Array_9_1_io_control_signal_mask = io_PE_control_1_mask; // @[PEArray.scala 274:40]
  assign PE_Array_9_2_clock = clock;
  assign PE_Array_9_2_reset = reset;
  assign PE_Array_9_2_io_FromAbovePE = PE_Array_9_1_io_ToBelowPE; // @[PEArray.scala 291:39]
  assign PE_Array_9_2_io_FromLeftPE = PE_Array_8_2_io_ToRightPE; // @[PEArray.scala 281:38]
  assign PE_Array_9_2_io_FromL1 = io_From_above_9; // @[PEArray.scala 308:32]
  assign PE_Array_9_2_io_control_signal_control = io_PE_control_2_control; // @[PEArray.scala 274:40]
  assign PE_Array_9_2_io_control_signal_count = io_PE_control_2_count; // @[PEArray.scala 274:40]
  assign PE_Array_9_2_io_control_signal_L0index = io_PE_control_2_L0index; // @[PEArray.scala 274:40]
  assign PE_Array_9_2_io_control_signal_mask = io_PE_control_2_mask; // @[PEArray.scala 274:40]
  assign PE_Array_9_2_io_control_signal_gru_out_width = io_PE_control_2_gru_out_width; // @[PEArray.scala 274:40]
  assign PE_Array_10_0_clock = clock;
  assign PE_Array_10_0_reset = reset;
  assign PE_Array_10_0_io_FromAbovePE = PE_Array_10_2_io_ToBelowPE; // @[PEArray.scala 297:35]
  assign PE_Array_10_0_io_FromLeftPE = PE_Array_9_0_io_ToRightPE; // @[PEArray.scala 281:38]
  assign PE_Array_10_0_io_FromL1 = io_From_above_10; // @[PEArray.scala 308:32]
  assign PE_Array_10_0_io_control_signal_mask = io_PE_control_0_mask; // @[PEArray.scala 274:40]
  assign PE_Array_10_1_clock = clock;
  assign PE_Array_10_1_reset = reset;
  assign PE_Array_10_1_io_FromAbovePE = PE_Array_10_0_io_ToBelowPE; // @[PEArray.scala 291:39]
  assign PE_Array_10_1_io_FromLeftPE = PE_Array_9_1_io_ToRightPE; // @[PEArray.scala 281:38]
  assign PE_Array_10_1_io_FromL1 = io_From_above_10; // @[PEArray.scala 308:32]
  assign PE_Array_10_1_io_control_signal_mask = io_PE_control_1_mask; // @[PEArray.scala 274:40]
  assign PE_Array_10_2_clock = clock;
  assign PE_Array_10_2_reset = reset;
  assign PE_Array_10_2_io_FromAbovePE = PE_Array_10_1_io_ToBelowPE; // @[PEArray.scala 291:39]
  assign PE_Array_10_2_io_FromLeftPE = PE_Array_9_2_io_ToRightPE; // @[PEArray.scala 281:38]
  assign PE_Array_10_2_io_FromL1 = io_From_above_10; // @[PEArray.scala 308:32]
  assign PE_Array_10_2_io_control_signal_control = io_PE_control_2_control; // @[PEArray.scala 274:40]
  assign PE_Array_10_2_io_control_signal_count = io_PE_control_2_count; // @[PEArray.scala 274:40]
  assign PE_Array_10_2_io_control_signal_L0index = io_PE_control_2_L0index; // @[PEArray.scala 274:40]
  assign PE_Array_10_2_io_control_signal_mask = io_PE_control_2_mask; // @[PEArray.scala 274:40]
  assign PE_Array_10_2_io_control_signal_gru_out_width = io_PE_control_2_gru_out_width; // @[PEArray.scala 274:40]
  assign PE_Array_11_0_clock = clock;
  assign PE_Array_11_0_reset = reset;
  assign PE_Array_11_0_io_FromAbovePE = PE_Array_11_2_io_ToBelowPE; // @[PEArray.scala 297:35]
  assign PE_Array_11_0_io_FromLeftPE = PE_Array_10_0_io_ToRightPE; // @[PEArray.scala 281:38]
  assign PE_Array_11_0_io_FromL1 = io_From_above_11; // @[PEArray.scala 308:32]
  assign PE_Array_11_0_io_control_signal_mask = io_PE_control_0_mask; // @[PEArray.scala 274:40]
  assign PE_Array_11_1_clock = clock;
  assign PE_Array_11_1_reset = reset;
  assign PE_Array_11_1_io_FromAbovePE = PE_Array_11_0_io_ToBelowPE; // @[PEArray.scala 291:39]
  assign PE_Array_11_1_io_FromLeftPE = PE_Array_10_1_io_ToRightPE; // @[PEArray.scala 281:38]
  assign PE_Array_11_1_io_FromL1 = io_From_above_11; // @[PEArray.scala 308:32]
  assign PE_Array_11_1_io_control_signal_mask = io_PE_control_1_mask; // @[PEArray.scala 274:40]
  assign PE_Array_11_2_clock = clock;
  assign PE_Array_11_2_reset = reset;
  assign PE_Array_11_2_io_FromAbovePE = PE_Array_11_1_io_ToBelowPE; // @[PEArray.scala 291:39]
  assign PE_Array_11_2_io_FromLeftPE = PE_Array_10_2_io_ToRightPE; // @[PEArray.scala 281:38]
  assign PE_Array_11_2_io_FromL1 = io_From_above_11; // @[PEArray.scala 308:32]
  assign PE_Array_11_2_io_control_signal_control = io_PE_control_2_control; // @[PEArray.scala 274:40]
  assign PE_Array_11_2_io_control_signal_count = io_PE_control_2_count; // @[PEArray.scala 274:40]
  assign PE_Array_11_2_io_control_signal_L0index = io_PE_control_2_L0index; // @[PEArray.scala 274:40]
  assign PE_Array_11_2_io_control_signal_mask = io_PE_control_2_mask; // @[PEArray.scala 274:40]
  assign PE_Array_11_2_io_control_signal_gru_out_width = io_PE_control_2_gru_out_width; // @[PEArray.scala 274:40]
  always @(posedge clock) begin
    rd_data_mux_delay <= io_rd_data_mux; // @[PEArray.scala 304:34]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rd_data_mux_delay = _RAND_0[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FSM(
  input         clock,
  input         reset,
  input         io_Start,
  input  [15:0] io_Input_Data,
  input         io_Input_Valid,
  output        io_Input_Ready,
  output [15:0] io_L1_wr_data,
  output        io_To_L1_control,
  output [11:0] io_L1_rd_addr_0,
  output [11:0] io_L1_rd_addr_1,
  output [11:0] io_L1_rd_addr_2,
  output [11:0] io_L1_rd_addr_3,
  output [11:0] io_L1_rd_addr_4,
  output [11:0] io_L1_rd_addr_5,
  output [11:0] io_L1_rd_addr_6,
  output [11:0] io_L1_rd_addr_7,
  output [11:0] io_L1_rd_addr_8,
  output [11:0] io_L1_rd_addr_9,
  output [11:0] io_L1_rd_addr_10,
  output [11:0] io_L1_rd_addr_11,
  output [3:0]  io_PE_rd_data_mux,
  output [11:0] io_L1_wr_addr_0,
  output [11:0] io_L1_wr_addr_1,
  output [11:0] io_L1_wr_addr_2,
  output [11:0] io_L1_wr_addr_3,
  output [11:0] io_L1_wr_addr_4,
  output [11:0] io_L1_wr_addr_5,
  output [11:0] io_L1_wr_addr_6,
  output [11:0] io_L1_wr_addr_7,
  output [11:0] io_L1_wr_addr_8,
  output [11:0] io_L1_wr_addr_9,
  output [11:0] io_L1_wr_addr_10,
  output [11:0] io_L1_wr_addr_11,
  output        io_L1_wrEna_0,
  output        io_L1_wrEna_1,
  output        io_L1_wrEna_2,
  output        io_L1_wrEna_3,
  output        io_L1_wrEna_4,
  output        io_L1_wrEna_5,
  output        io_L1_wrEna_6,
  output        io_L1_wrEna_7,
  output        io_L1_wrEna_8,
  output        io_L1_wrEna_9,
  output        io_L1_wrEna_10,
  output        io_L1_wrEna_11,
  output [11:0] io_PEArray_ctrl_0_mask,
  output [11:0] io_PEArray_ctrl_1_mask,
  output [2:0]  io_PEArray_ctrl_2_control,
  output [9:0]  io_PEArray_ctrl_2_count,
  output [5:0]  io_PEArray_ctrl_2_L0index,
  output [11:0] io_PEArray_ctrl_2_mask,
  output [7:0]  io_PEArray_ctrl_2_gru_out_width,
  output [1:0]  io_BNArray_ctrl_0,
  output [1:0]  io_BNArray_ctrl_1,
  output [1:0]  io_BNArray_ctrl_2,
  output [1:0]  io_BNArray_ctrl_3,
  output [1:0]  io_BNArray_ctrl_4,
  output [1:0]  io_BNArray_ctrl_5,
  output [1:0]  io_BNArray_ctrl_6,
  output [1:0]  io_BNArray_ctrl_7,
  output [1:0]  io_BNArray_ctrl_8,
  output [1:0]  io_BNArray_ctrl_9,
  output [1:0]  io_BNArray_ctrl_10,
  output [1:0]  io_BNArray_ctrl_11,
  output [1:0]  io_BN_Unit_ctrl,
  output        io_Relu6Array_ctrl_0,
  output        io_Relu6Array_ctrl_1,
  output        io_Relu6Array_ctrl_2,
  output        io_Relu6Array_ctrl_3,
  output        io_Relu6Array_ctrl_4,
  output        io_Relu6Array_ctrl_5,
  output        io_Relu6Array_ctrl_6,
  output        io_Relu6Array_ctrl_7,
  output        io_Relu6Array_ctrl_8,
  output        io_Relu6Array_ctrl_9,
  output        io_Relu6Array_ctrl_10,
  output        io_Relu6Array_ctrl_11,
  output [1:0]  io_PE_above_data_ctrl,
  output [1:0]  io_Activation_ctrl,
  output [2:0]  io_Ht_to_PE_control,
  output        io_Ht_wrEna,
  output [5:0]  io_Ht_wrAddr,
  output [5:0]  io_Zt_rdAddr,
  output        io_Zt_wrEna,
  output [5:0]  io_Zt_wrAddr,
  output [5:0]  io_Rt_rdAddr,
  output        io_Rt_wrEna,
  output [5:0]  io_Rt_wrAddr,
  output [5:0]  io_WhXt_rdAddr,
  output        io_WhXt_wrEna,
  output [5:0]  io_WhXt_wrAddr,
  output [5:0]  io_Uhht_1_rdAddr,
  output        io_Uhht_1_wrEna,
  output [5:0]  io_Uhht_1_wrAddr,
  output [2:0]  io_FC_temp_to_PE_control,
  output        io_FC_temp_wrEna,
  output [5:0]  io_FC_temp_wrAddr,
  output        io_Result_wrEna,
  output [3:0]  io_Result_wrAddr
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
`endif // RANDOMIZE_REG_INIT
  reg [11:0] L1_rd_addr_0; // @[FSM.scala 60:28]
  reg [11:0] L1_rd_addr_1; // @[FSM.scala 60:28]
  reg [11:0] L1_rd_addr_2; // @[FSM.scala 60:28]
  reg [11:0] L1_rd_addr_3; // @[FSM.scala 60:28]
  reg [11:0] L1_rd_addr_4; // @[FSM.scala 60:28]
  reg [11:0] L1_rd_addr_5; // @[FSM.scala 60:28]
  reg [11:0] L1_rd_addr_6; // @[FSM.scala 60:28]
  reg [11:0] L1_rd_addr_7; // @[FSM.scala 60:28]
  reg [11:0] L1_rd_addr_8; // @[FSM.scala 60:28]
  reg [11:0] L1_rd_addr_9; // @[FSM.scala 60:28]
  reg [11:0] L1_rd_addr_10; // @[FSM.scala 60:28]
  reg [11:0] L1_rd_addr_11; // @[FSM.scala 60:28]
  reg [3:0] PE_rd_data_mux; // @[FSM.scala 61:32]
  reg [11:0] L1_wr_addr_0; // @[FSM.scala 62:28]
  reg [11:0] L1_wr_addr_1; // @[FSM.scala 62:28]
  reg [11:0] L1_wr_addr_2; // @[FSM.scala 62:28]
  reg [11:0] L1_wr_addr_3; // @[FSM.scala 62:28]
  reg [11:0] L1_wr_addr_4; // @[FSM.scala 62:28]
  reg [11:0] L1_wr_addr_5; // @[FSM.scala 62:28]
  reg [11:0] L1_wr_addr_6; // @[FSM.scala 62:28]
  reg [11:0] L1_wr_addr_7; // @[FSM.scala 62:28]
  reg [11:0] L1_wr_addr_8; // @[FSM.scala 62:28]
  reg [11:0] L1_wr_addr_9; // @[FSM.scala 62:28]
  reg [11:0] L1_wr_addr_10; // @[FSM.scala 62:28]
  reg [11:0] L1_wr_addr_11; // @[FSM.scala 62:28]
  reg  L1_wrEna_0; // @[FSM.scala 63:28]
  reg  L1_wrEna_1; // @[FSM.scala 63:28]
  reg  L1_wrEna_2; // @[FSM.scala 63:28]
  reg  L1_wrEna_3; // @[FSM.scala 63:28]
  reg  L1_wrEna_4; // @[FSM.scala 63:28]
  reg  L1_wrEna_5; // @[FSM.scala 63:28]
  reg  L1_wrEna_6; // @[FSM.scala 63:28]
  reg  L1_wrEna_7; // @[FSM.scala 63:28]
  reg  L1_wrEna_8; // @[FSM.scala 63:28]
  reg  L1_wrEna_9; // @[FSM.scala 63:28]
  reg  L1_wrEna_10; // @[FSM.scala 63:28]
  reg  L1_wrEna_11; // @[FSM.scala 63:28]
  reg [11:0] PEArray_ctrl_0_mask; // @[FSM.scala 64:28]
  reg [11:0] PEArray_ctrl_1_mask; // @[FSM.scala 64:28]
  reg [2:0] PEArray_ctrl_2_control; // @[FSM.scala 64:28]
  reg [9:0] PEArray_ctrl_2_count; // @[FSM.scala 64:28]
  reg [5:0] PEArray_ctrl_2_L0index; // @[FSM.scala 64:28]
  reg [11:0] PEArray_ctrl_2_mask; // @[FSM.scala 64:28]
  reg [7:0] PEArray_ctrl_2_gru_out_width; // @[FSM.scala 64:28]
  reg [1:0] BNArray_ctrl_0; // @[FSM.scala 65:28]
  reg [1:0] BNArray_ctrl_1; // @[FSM.scala 65:28]
  reg [1:0] BNArray_ctrl_2; // @[FSM.scala 65:28]
  reg [1:0] BNArray_ctrl_3; // @[FSM.scala 65:28]
  reg [1:0] BNArray_ctrl_4; // @[FSM.scala 65:28]
  reg [1:0] BNArray_ctrl_5; // @[FSM.scala 65:28]
  reg [1:0] BNArray_ctrl_6; // @[FSM.scala 65:28]
  reg [1:0] BNArray_ctrl_7; // @[FSM.scala 65:28]
  reg [1:0] BNArray_ctrl_8; // @[FSM.scala 65:28]
  reg [1:0] BNArray_ctrl_9; // @[FSM.scala 65:28]
  reg [1:0] BNArray_ctrl_10; // @[FSM.scala 65:28]
  reg [1:0] BNArray_ctrl_11; // @[FSM.scala 65:28]
  reg [1:0] BN_Unit_ctrl; // @[FSM.scala 69:28]
  reg  Relu6Array_ctrl_0; // @[FSM.scala 73:28]
  reg  Relu6Array_ctrl_1; // @[FSM.scala 73:28]
  reg  Relu6Array_ctrl_2; // @[FSM.scala 73:28]
  reg  Relu6Array_ctrl_3; // @[FSM.scala 73:28]
  reg  Relu6Array_ctrl_4; // @[FSM.scala 73:28]
  reg  Relu6Array_ctrl_5; // @[FSM.scala 73:28]
  reg  Relu6Array_ctrl_6; // @[FSM.scala 73:28]
  reg  Relu6Array_ctrl_7; // @[FSM.scala 73:28]
  reg  Relu6Array_ctrl_8; // @[FSM.scala 73:28]
  reg  Relu6Array_ctrl_9; // @[FSM.scala 73:28]
  reg  Relu6Array_ctrl_10; // @[FSM.scala 73:28]
  reg  Relu6Array_ctrl_11; // @[FSM.scala 73:28]
  reg [1:0] PE_above_data_ctrl; // @[FSM.scala 74:35]
  reg [1:0] Activation_ctrl; // @[FSM.scala 75:32]
  reg [2:0] Ht_to_PE_control; // @[FSM.scala 77:36]
  reg  Ht_wrEna; // @[FSM.scala 79:36]
  reg [5:0] Ht_wrAddr; // @[FSM.scala 80:36]
  reg [5:0] Zt_rdAddr; // @[FSM.scala 81:36]
  reg  Zt_wrEna; // @[FSM.scala 82:36]
  reg [5:0] Zt_wrAddr; // @[FSM.scala 83:36]
  reg [5:0] Rt_rdAddr; // @[FSM.scala 84:36]
  reg  Rt_wrEna; // @[FSM.scala 85:36]
  reg [5:0] Rt_wrAddr; // @[FSM.scala 86:36]
  reg [5:0] WhXt_rdAddr; // @[FSM.scala 87:36]
  reg  WhXt_wrEna; // @[FSM.scala 88:36]
  reg [5:0] WhXt_wrAddr; // @[FSM.scala 89:36]
  reg [5:0] Uhht_1_rdAddr; // @[FSM.scala 90:36]
  reg  Uhht_1_wrEna; // @[FSM.scala 91:36]
  reg [5:0] Uhht_1_wrAddr; // @[FSM.scala 92:36]
  reg [2:0] FC_temp_to_PE_control; // @[FSM.scala 94:38]
  reg  FC_temp_wrEna; // @[FSM.scala 96:38]
  reg [5:0] FC_temp_wrAddr; // @[FSM.scala 97:38]
  reg  Result_wrEna; // @[FSM.scala 99:38]
  reg [3:0] Result_wrAddr; // @[FSM.scala 100:38]
  reg [15:0] Data_temp; // @[FSM.scala 104:22]
  reg  Data_temp_used; // @[FSM.scala 105:31]
  reg [15:0] L1_wr_data; // @[FSM.scala 106:27]
  reg [2:0] state; // @[FSM.scala 159:22]
  reg [3:0] gru_state; // @[FSM.scala 160:26]
  reg [9:0] count; // @[FSM.scala 161:22]
  reg [6:0] count1; // @[FSM.scala 162:23]
  reg [5:0] gru_count; // @[FSM.scala 164:26]
  reg [3:0] read_index; // @[FSM.scala 165:27]
  reg [1:0] fc_state; // @[FSM.scala 166:25]
  wire  _T = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_2 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_3 = count == 10'h0; // @[FSM.scala 175:18]
  wire  _T_5 = count == 10'h1; // @[FSM.scala 182:20]
  wire [15:0] _GEN_3 = count == 10'h1 ? Data_temp : L1_wr_data; // @[FSM.scala 182:28 FSM.scala 183:22 FSM.scala 106:27]
  wire [11:0] _GEN_4 = count == 10'h1 ? 12'h1b8 : L1_wr_addr_0; // @[FSM.scala 182:28 FSM.scala 185:27 FSM.scala 62:28]
  wire  _GEN_5 = count == 10'h1 | L1_wrEna_0; // @[FSM.scala 182:28 FSM.scala 186:25 FSM.scala 63:28]
  wire [11:0] _GEN_6 = count == 10'h1 ? 12'h1b8 : L1_wr_addr_1; // @[FSM.scala 182:28 FSM.scala 185:27 FSM.scala 62:28]
  wire  _GEN_7 = count == 10'h1 | L1_wrEna_1; // @[FSM.scala 182:28 FSM.scala 186:25 FSM.scala 63:28]
  wire [11:0] _GEN_8 = count == 10'h1 ? 12'h1b8 : L1_wr_addr_2; // @[FSM.scala 182:28 FSM.scala 185:27 FSM.scala 62:28]
  wire  _GEN_9 = count == 10'h1 | L1_wrEna_2; // @[FSM.scala 182:28 FSM.scala 186:25 FSM.scala 63:28]
  wire [11:0] _GEN_10 = count == 10'h1 ? 12'h1b8 : L1_wr_addr_3; // @[FSM.scala 182:28 FSM.scala 185:27 FSM.scala 62:28]
  wire  _GEN_11 = count == 10'h1 | L1_wrEna_3; // @[FSM.scala 182:28 FSM.scala 186:25 FSM.scala 63:28]
  wire [11:0] _GEN_12 = count == 10'h1 ? 12'h1b8 : L1_wr_addr_4; // @[FSM.scala 182:28 FSM.scala 185:27 FSM.scala 62:28]
  wire  _GEN_13 = count == 10'h1 | L1_wrEna_4; // @[FSM.scala 182:28 FSM.scala 186:25 FSM.scala 63:28]
  wire [11:0] _GEN_14 = count == 10'h1 ? 12'h1b8 : L1_wr_addr_5; // @[FSM.scala 182:28 FSM.scala 185:27 FSM.scala 62:28]
  wire  _GEN_15 = count == 10'h1 | L1_wrEna_5; // @[FSM.scala 182:28 FSM.scala 186:25 FSM.scala 63:28]
  wire [11:0] _GEN_16 = count == 10'h1 ? 12'h1b8 : L1_wr_addr_6; // @[FSM.scala 182:28 FSM.scala 185:27 FSM.scala 62:28]
  wire  _GEN_17 = count == 10'h1 | L1_wrEna_6; // @[FSM.scala 182:28 FSM.scala 186:25 FSM.scala 63:28]
  wire [11:0] _GEN_18 = count == 10'h1 ? 12'h1b8 : L1_wr_addr_7; // @[FSM.scala 182:28 FSM.scala 185:27 FSM.scala 62:28]
  wire  _GEN_19 = count == 10'h1 | L1_wrEna_7; // @[FSM.scala 182:28 FSM.scala 186:25 FSM.scala 63:28]
  wire [11:0] _GEN_20 = count == 10'h1 ? 12'h1b8 : L1_wr_addr_8; // @[FSM.scala 182:28 FSM.scala 185:27 FSM.scala 62:28]
  wire  _GEN_21 = count == 10'h1 | L1_wrEna_8; // @[FSM.scala 182:28 FSM.scala 186:25 FSM.scala 63:28]
  wire [11:0] _GEN_22 = count == 10'h1 ? 12'h1b8 : L1_wr_addr_9; // @[FSM.scala 182:28 FSM.scala 185:27 FSM.scala 62:28]
  wire  _GEN_23 = count == 10'h1 | L1_wrEna_9; // @[FSM.scala 182:28 FSM.scala 186:25 FSM.scala 63:28]
  wire [11:0] _GEN_24 = count == 10'h1 ? 12'h1b8 : L1_wr_addr_10; // @[FSM.scala 182:28 FSM.scala 185:27 FSM.scala 62:28]
  wire  _GEN_25 = count == 10'h1 | L1_wrEna_10; // @[FSM.scala 182:28 FSM.scala 186:25 FSM.scala 63:28]
  wire [11:0] _GEN_26 = count == 10'h1 ? 12'h1b8 : L1_wr_addr_11; // @[FSM.scala 182:28 FSM.scala 185:27 FSM.scala 62:28]
  wire  _GEN_27 = count == 10'h1 | L1_wrEna_11; // @[FSM.scala 182:28 FSM.scala 186:25 FSM.scala 63:28]
  wire [11:0] _L1_wr_addr_0_T_1 = L1_wr_addr_0 + 12'h1; // @[FSM.scala 192:44]
  wire [11:0] _L1_wr_addr_1_T_1 = L1_wr_addr_1 + 12'h1; // @[FSM.scala 192:44]
  wire [11:0] _L1_wr_addr_2_T_1 = L1_wr_addr_2 + 12'h1; // @[FSM.scala 192:44]
  wire [11:0] _L1_wr_addr_3_T_1 = L1_wr_addr_3 + 12'h1; // @[FSM.scala 192:44]
  wire [11:0] _L1_wr_addr_4_T_1 = L1_wr_addr_4 + 12'h1; // @[FSM.scala 192:44]
  wire [11:0] _L1_wr_addr_5_T_1 = L1_wr_addr_5 + 12'h1; // @[FSM.scala 192:44]
  wire [11:0] _L1_wr_addr_6_T_1 = L1_wr_addr_6 + 12'h1; // @[FSM.scala 192:44]
  wire [11:0] _L1_wr_addr_7_T_1 = L1_wr_addr_7 + 12'h1; // @[FSM.scala 192:44]
  wire [11:0] _L1_wr_addr_8_T_1 = L1_wr_addr_8 + 12'h1; // @[FSM.scala 192:44]
  wire [11:0] _L1_wr_addr_9_T_1 = L1_wr_addr_9 + 12'h1; // @[FSM.scala 192:44]
  wire [11:0] _L1_wr_addr_10_T_1 = L1_wr_addr_10 + 12'h1; // @[FSM.scala 192:44]
  wire [11:0] _L1_wr_addr_11_T_1 = L1_wr_addr_11 + 12'h1; // @[FSM.scala 192:44]
  wire  _GEN_30 = count >= 10'h2 & count <= 10'hf | _GEN_5; // @[FSM.scala 189:44 FSM.scala 193:25]
  wire  _GEN_32 = count >= 10'h2 & count <= 10'hf | _GEN_7; // @[FSM.scala 189:44 FSM.scala 193:25]
  wire  _GEN_34 = count >= 10'h2 & count <= 10'hf | _GEN_9; // @[FSM.scala 189:44 FSM.scala 193:25]
  wire  _GEN_36 = count >= 10'h2 & count <= 10'hf | _GEN_11; // @[FSM.scala 189:44 FSM.scala 193:25]
  wire  _GEN_38 = count >= 10'h2 & count <= 10'hf | _GEN_13; // @[FSM.scala 189:44 FSM.scala 193:25]
  wire  _GEN_40 = count >= 10'h2 & count <= 10'hf | _GEN_15; // @[FSM.scala 189:44 FSM.scala 193:25]
  wire  _GEN_42 = count >= 10'h2 & count <= 10'hf | _GEN_17; // @[FSM.scala 189:44 FSM.scala 193:25]
  wire  _GEN_44 = count >= 10'h2 & count <= 10'hf | _GEN_19; // @[FSM.scala 189:44 FSM.scala 193:25]
  wire  _GEN_46 = count >= 10'h2 & count <= 10'hf | _GEN_21; // @[FSM.scala 189:44 FSM.scala 193:25]
  wire  _GEN_48 = count >= 10'h2 & count <= 10'hf | _GEN_23; // @[FSM.scala 189:44 FSM.scala 193:25]
  wire  _GEN_50 = count >= 10'h2 & count <= 10'hf | _GEN_25; // @[FSM.scala 189:44 FSM.scala 193:25]
  wire  _GEN_52 = count >= 10'h2 & count <= 10'hf | _GEN_27; // @[FSM.scala 189:44 FSM.scala 193:25]
  wire  _GEN_53 = ~Data_temp_used | Data_temp_used; // @[FSM.scala 179:39 FSM.scala 180:24 FSM.scala 105:31]
  wire  _GEN_56 = ~Data_temp_used & _GEN_30; // @[FSM.scala 179:39 FSM.scala 198:23]
  wire  _GEN_58 = ~Data_temp_used & _GEN_32; // @[FSM.scala 179:39 FSM.scala 198:23]
  wire  _GEN_60 = ~Data_temp_used & _GEN_34; // @[FSM.scala 179:39 FSM.scala 198:23]
  wire  _GEN_62 = ~Data_temp_used & _GEN_36; // @[FSM.scala 179:39 FSM.scala 198:23]
  wire  _GEN_64 = ~Data_temp_used & _GEN_38; // @[FSM.scala 179:39 FSM.scala 198:23]
  wire  _GEN_66 = ~Data_temp_used & _GEN_40; // @[FSM.scala 179:39 FSM.scala 198:23]
  wire  _GEN_68 = ~Data_temp_used & _GEN_42; // @[FSM.scala 179:39 FSM.scala 198:23]
  wire  _GEN_70 = ~Data_temp_used & _GEN_44; // @[FSM.scala 179:39 FSM.scala 198:23]
  wire  _GEN_72 = ~Data_temp_used & _GEN_46; // @[FSM.scala 179:39 FSM.scala 198:23]
  wire  _GEN_74 = ~Data_temp_used & _GEN_48; // @[FSM.scala 179:39 FSM.scala 198:23]
  wire  _GEN_76 = ~Data_temp_used & _GEN_50; // @[FSM.scala 179:39 FSM.scala 198:23]
  wire  _GEN_78 = ~Data_temp_used & _GEN_52; // @[FSM.scala 179:39 FSM.scala 198:23]
  wire [9:0] _count_T_1 = count + 10'h1; // @[FSM.scala 205:24]
  wire  _GEN_80 = io_Input_Valid & io_Input_Ready ? 1'h0 : _GEN_53; // @[FSM.scala 202:67 FSM.scala 204:24]
  wire  _GEN_83 = count == 10'h10 ? 1'h0 : _T_3; // @[FSM.scala 207:27 FSM.scala 209:26]
  wire  _T_13 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire [9:0] _GEN_84 = count != 10'h34 ? _count_T_1 : count; // @[FSM.scala 214:27 FSM.scala 215:15 FSM.scala 161:22]
  wire [6:0] _count1_T_1 = count1 + 7'h1; // @[FSM.scala 218:26]
  wire [6:0] _GEN_85 = count1 != 7'h9 ? _count1_T_1 : 7'h0; // @[FSM.scala 217:27 FSM.scala 218:16 FSM.scala 220:16]
  wire [11:0] _GEN_87 = _T_3 ? 12'hfff : PEArray_ctrl_0_mask; // @[FSM.scala 223:26 FSM.scala 226:32 FSM.scala 64:28]
  wire [11:0] _GEN_89 = _T_3 ? 12'hfff : PEArray_ctrl_1_mask; // @[FSM.scala 223:26 FSM.scala 226:32 FSM.scala 64:28]
  wire [11:0] _GEN_91 = _T_3 ? 12'hfff : PEArray_ctrl_2_mask; // @[FSM.scala 223:26 FSM.scala 226:32 FSM.scala 64:28]
  wire [11:0] _GEN_92 = _T_3 ? 12'h0 : L1_rd_addr_0; // @[FSM.scala 223:26 FSM.scala 230:25 FSM.scala 60:28]
  wire [11:0] _GEN_93 = _T_3 ? 12'h0 : L1_rd_addr_1; // @[FSM.scala 223:26 FSM.scala 230:25 FSM.scala 60:28]
  wire [11:0] _GEN_94 = _T_3 ? 12'h0 : L1_rd_addr_2; // @[FSM.scala 223:26 FSM.scala 230:25 FSM.scala 60:28]
  wire [11:0] _GEN_95 = _T_3 ? 12'h0 : L1_rd_addr_3; // @[FSM.scala 223:26 FSM.scala 230:25 FSM.scala 60:28]
  wire [11:0] _GEN_96 = _T_3 ? 12'h0 : L1_rd_addr_4; // @[FSM.scala 223:26 FSM.scala 230:25 FSM.scala 60:28]
  wire [11:0] _GEN_97 = _T_3 ? 12'h0 : L1_rd_addr_5; // @[FSM.scala 223:26 FSM.scala 230:25 FSM.scala 60:28]
  wire [11:0] _GEN_98 = _T_3 ? 12'h0 : L1_rd_addr_6; // @[FSM.scala 223:26 FSM.scala 230:25 FSM.scala 60:28]
  wire [11:0] _GEN_99 = _T_3 ? 12'h0 : L1_rd_addr_7; // @[FSM.scala 223:26 FSM.scala 230:25 FSM.scala 60:28]
  wire [11:0] _GEN_100 = _T_3 ? 12'h0 : L1_rd_addr_8; // @[FSM.scala 223:26 FSM.scala 230:25 FSM.scala 60:28]
  wire [11:0] _GEN_101 = _T_3 ? 12'h0 : L1_rd_addr_9; // @[FSM.scala 223:26 FSM.scala 230:25 FSM.scala 60:28]
  wire [11:0] _GEN_102 = _T_3 ? 12'h0 : L1_rd_addr_10; // @[FSM.scala 223:26 FSM.scala 230:25 FSM.scala 60:28]
  wire [11:0] _GEN_103 = _T_3 ? 12'h0 : L1_rd_addr_11; // @[FSM.scala 223:26 FSM.scala 230:25 FSM.scala 60:28]
  wire [1:0] _GEN_104 = _T_3 ? 2'h0 : PE_above_data_ctrl; // @[FSM.scala 223:26 FSM.scala 232:28 FSM.scala 74:35]
  wire [3:0] _GEN_105 = _T_3 ? 4'h0 : PE_rd_data_mux; // @[FSM.scala 223:26 FSM.scala 233:24 FSM.scala 61:32]
  wire [11:0] _GEN_108 = _T_5 ? 12'h0 : _GEN_91; // @[FSM.scala 235:26 FSM.scala 237:32]
  wire  _T_18 = count >= 10'h1; // @[FSM.scala 241:19]
  wire [11:0] _L1_rd_addr_0_T_1 = L1_rd_addr_0 + 12'h1; // @[FSM.scala 243:42]
  wire [11:0] _L1_rd_addr_1_T_1 = L1_rd_addr_1 + 12'h1; // @[FSM.scala 243:42]
  wire [11:0] _L1_rd_addr_2_T_1 = L1_rd_addr_2 + 12'h1; // @[FSM.scala 243:42]
  wire [11:0] _L1_rd_addr_3_T_1 = L1_rd_addr_3 + 12'h1; // @[FSM.scala 243:42]
  wire [11:0] _L1_rd_addr_4_T_1 = L1_rd_addr_4 + 12'h1; // @[FSM.scala 243:42]
  wire [11:0] _L1_rd_addr_5_T_1 = L1_rd_addr_5 + 12'h1; // @[FSM.scala 243:42]
  wire [11:0] _L1_rd_addr_6_T_1 = L1_rd_addr_6 + 12'h1; // @[FSM.scala 243:42]
  wire [11:0] _L1_rd_addr_7_T_1 = L1_rd_addr_7 + 12'h1; // @[FSM.scala 243:42]
  wire [11:0] _L1_rd_addr_8_T_1 = L1_rd_addr_8 + 12'h1; // @[FSM.scala 243:42]
  wire [11:0] _L1_rd_addr_9_T_1 = L1_rd_addr_9 + 12'h1; // @[FSM.scala 243:42]
  wire [11:0] _L1_rd_addr_10_T_1 = L1_rd_addr_10 + 12'h1; // @[FSM.scala 243:42]
  wire [11:0] _L1_rd_addr_11_T_1 = L1_rd_addr_11 + 12'h1; // @[FSM.scala 243:42]
  wire  _T_21 = count == 10'h4; // @[FSM.scala 247:18]
  wire  _GEN_121 = count == 10'h4 | L1_wrEna_0; // @[FSM.scala 247:26 FSM.scala 249:23 FSM.scala 63:28]
  wire [11:0] _GEN_122 = count == 10'h4 ? 12'h190 : L1_wr_addr_0; // @[FSM.scala 247:26 FSM.scala 250:25 FSM.scala 62:28]
  wire  _GEN_125 = count == 10'h4 | L1_wrEna_1; // @[FSM.scala 247:26 FSM.scala 249:23 FSM.scala 63:28]
  wire [11:0] _GEN_126 = count == 10'h4 ? 12'h190 : L1_wr_addr_1; // @[FSM.scala 247:26 FSM.scala 250:25 FSM.scala 62:28]
  wire  _GEN_129 = count == 10'h4 | L1_wrEna_2; // @[FSM.scala 247:26 FSM.scala 249:23 FSM.scala 63:28]
  wire [11:0] _GEN_130 = count == 10'h4 ? 12'h190 : L1_wr_addr_2; // @[FSM.scala 247:26 FSM.scala 250:25 FSM.scala 62:28]
  wire  _GEN_133 = count == 10'h4 | L1_wrEna_3; // @[FSM.scala 247:26 FSM.scala 249:23 FSM.scala 63:28]
  wire [11:0] _GEN_134 = count == 10'h4 ? 12'h190 : L1_wr_addr_3; // @[FSM.scala 247:26 FSM.scala 250:25 FSM.scala 62:28]
  wire  _GEN_137 = count == 10'h4 | L1_wrEna_4; // @[FSM.scala 247:26 FSM.scala 249:23 FSM.scala 63:28]
  wire [11:0] _GEN_138 = count == 10'h4 ? 12'h190 : L1_wr_addr_4; // @[FSM.scala 247:26 FSM.scala 250:25 FSM.scala 62:28]
  wire  _GEN_141 = count == 10'h4 | L1_wrEna_5; // @[FSM.scala 247:26 FSM.scala 249:23 FSM.scala 63:28]
  wire [11:0] _GEN_142 = count == 10'h4 ? 12'h190 : L1_wr_addr_5; // @[FSM.scala 247:26 FSM.scala 250:25 FSM.scala 62:28]
  wire  _GEN_145 = count == 10'h4 | L1_wrEna_6; // @[FSM.scala 247:26 FSM.scala 249:23 FSM.scala 63:28]
  wire [11:0] _GEN_146 = count == 10'h4 ? 12'h190 : L1_wr_addr_6; // @[FSM.scala 247:26 FSM.scala 250:25 FSM.scala 62:28]
  wire  _GEN_149 = count == 10'h4 | L1_wrEna_7; // @[FSM.scala 247:26 FSM.scala 249:23 FSM.scala 63:28]
  wire [11:0] _GEN_150 = count == 10'h4 ? 12'h190 : L1_wr_addr_7; // @[FSM.scala 247:26 FSM.scala 250:25 FSM.scala 62:28]
  wire  _GEN_153 = count == 10'h4 | L1_wrEna_8; // @[FSM.scala 247:26 FSM.scala 249:23 FSM.scala 63:28]
  wire [11:0] _GEN_154 = count == 10'h4 ? 12'h190 : L1_wr_addr_8; // @[FSM.scala 247:26 FSM.scala 250:25 FSM.scala 62:28]
  wire  _GEN_157 = count == 10'h4 | L1_wrEna_9; // @[FSM.scala 247:26 FSM.scala 249:23 FSM.scala 63:28]
  wire [11:0] _GEN_158 = count == 10'h4 ? 12'h190 : L1_wr_addr_9; // @[FSM.scala 247:26 FSM.scala 250:25 FSM.scala 62:28]
  wire  _GEN_161 = count == 10'h4 | L1_wrEna_10; // @[FSM.scala 247:26 FSM.scala 249:23 FSM.scala 63:28]
  wire [11:0] _GEN_162 = count == 10'h4 ? 12'h190 : L1_wr_addr_10; // @[FSM.scala 247:26 FSM.scala 250:25 FSM.scala 62:28]
  wire  _GEN_165 = count == 10'h4 | L1_wrEna_11; // @[FSM.scala 247:26 FSM.scala 249:23 FSM.scala 63:28]
  wire [11:0] _GEN_166 = count == 10'h4 ? 12'h190 : L1_wr_addr_11; // @[FSM.scala 247:26 FSM.scala 250:25 FSM.scala 62:28]
  wire  _T_25 = count1 == 7'h2; // @[FSM.scala 257:22]
  wire  _GEN_169 = count1 == 7'h2 & count1 == 7'h3 ? 1'h0 : 1'h1; // @[FSM.scala 257:51 FSM.scala 259:25 FSM.scala 263:25]
  wire [11:0] _GEN_170 = count1 == 7'h2 & count1 == 7'h3 ? _GEN_122 : _L1_wr_addr_0_T_1; // @[FSM.scala 257:51 FSM.scala 264:27]
  wire [11:0] _GEN_171 = count1 == 7'h2 & count1 == 7'h3 ? _GEN_126 : _L1_wr_addr_1_T_1; // @[FSM.scala 257:51 FSM.scala 264:27]
  wire [11:0] _GEN_172 = count1 == 7'h2 & count1 == 7'h3 ? _GEN_130 : _L1_wr_addr_2_T_1; // @[FSM.scala 257:51 FSM.scala 264:27]
  wire [11:0] _GEN_173 = count1 == 7'h2 & count1 == 7'h3 ? _GEN_134 : _L1_wr_addr_3_T_1; // @[FSM.scala 257:51 FSM.scala 264:27]
  wire [11:0] _GEN_174 = count1 == 7'h2 & count1 == 7'h3 ? _GEN_138 : _L1_wr_addr_4_T_1; // @[FSM.scala 257:51 FSM.scala 264:27]
  wire [11:0] _GEN_175 = count1 == 7'h2 & count1 == 7'h3 ? _GEN_142 : _L1_wr_addr_5_T_1; // @[FSM.scala 257:51 FSM.scala 264:27]
  wire [11:0] _GEN_176 = count1 == 7'h2 & count1 == 7'h3 ? _GEN_146 : _L1_wr_addr_6_T_1; // @[FSM.scala 257:51 FSM.scala 264:27]
  wire [11:0] _GEN_177 = count1 == 7'h2 & count1 == 7'h3 ? _GEN_150 : _L1_wr_addr_7_T_1; // @[FSM.scala 257:51 FSM.scala 264:27]
  wire [11:0] _GEN_178 = count1 == 7'h2 & count1 == 7'h3 ? _GEN_154 : _L1_wr_addr_8_T_1; // @[FSM.scala 257:51 FSM.scala 264:27]
  wire [11:0] _GEN_179 = count1 == 7'h2 & count1 == 7'h3 ? _GEN_158 : _L1_wr_addr_9_T_1; // @[FSM.scala 257:51 FSM.scala 264:27]
  wire [11:0] _GEN_180 = count1 == 7'h2 & count1 == 7'h3 ? _GEN_162 : _L1_wr_addr_10_T_1; // @[FSM.scala 257:51 FSM.scala 264:27]
  wire [11:0] _GEN_181 = count1 == 7'h2 & count1 == 7'h3 ? _GEN_166 : _L1_wr_addr_11_T_1; // @[FSM.scala 257:51 FSM.scala 264:27]
  wire  _GEN_182 = count >= 10'h5 & count <= 10'h2b ? _GEN_169 : _GEN_121; // @[FSM.scala 256:46]
  wire  _GEN_183 = count >= 10'h5 & count <= 10'h2b ? _GEN_169 : _GEN_125; // @[FSM.scala 256:46]
  wire  _GEN_184 = count >= 10'h5 & count <= 10'h2b ? _GEN_169 : _GEN_129; // @[FSM.scala 256:46]
  wire  _GEN_185 = count >= 10'h5 & count <= 10'h2b ? _GEN_169 : _GEN_133; // @[FSM.scala 256:46]
  wire  _GEN_186 = count >= 10'h5 & count <= 10'h2b ? _GEN_169 : _GEN_137; // @[FSM.scala 256:46]
  wire  _GEN_187 = count >= 10'h5 & count <= 10'h2b ? _GEN_169 : _GEN_141; // @[FSM.scala 256:46]
  wire  _GEN_188 = count >= 10'h5 & count <= 10'h2b ? _GEN_169 : _GEN_145; // @[FSM.scala 256:46]
  wire  _GEN_189 = count >= 10'h5 & count <= 10'h2b ? _GEN_169 : _GEN_149; // @[FSM.scala 256:46]
  wire  _GEN_190 = count >= 10'h5 & count <= 10'h2b ? _GEN_169 : _GEN_153; // @[FSM.scala 256:46]
  wire  _GEN_191 = count >= 10'h5 & count <= 10'h2b ? _GEN_169 : _GEN_157; // @[FSM.scala 256:46]
  wire  _GEN_192 = count >= 10'h5 & count <= 10'h2b ? _GEN_169 : _GEN_161; // @[FSM.scala 256:46]
  wire  _GEN_193 = count >= 10'h5 & count <= 10'h2b ? _GEN_169 : _GEN_165; // @[FSM.scala 256:46]
  wire [11:0] _GEN_194 = count >= 10'h5 & count <= 10'h2b ? _GEN_170 : _GEN_122; // @[FSM.scala 256:46]
  wire  _GEN_206 = count >= 10'h2c & count <= 10'h33 | _GEN_182; // @[FSM.scala 268:47 FSM.scala 269:21]
  wire  _GEN_208 = count >= 10'h2c & count <= 10'h33 ? 1'h0 : _GEN_183; // @[FSM.scala 268:47 FSM.scala 272:23]
  wire  _GEN_209 = count >= 10'h2c & count <= 10'h33 ? 1'h0 : _GEN_184; // @[FSM.scala 268:47 FSM.scala 272:23]
  wire  _GEN_210 = count >= 10'h2c & count <= 10'h33 ? 1'h0 : _GEN_185; // @[FSM.scala 268:47 FSM.scala 272:23]
  wire  _GEN_211 = count >= 10'h2c & count <= 10'h33 ? 1'h0 : _GEN_186; // @[FSM.scala 268:47 FSM.scala 272:23]
  wire  _GEN_212 = count >= 10'h2c & count <= 10'h33 ? 1'h0 : _GEN_187; // @[FSM.scala 268:47 FSM.scala 272:23]
  wire  _GEN_213 = count >= 10'h2c & count <= 10'h33 ? 1'h0 : _GEN_188; // @[FSM.scala 268:47 FSM.scala 272:23]
  wire  _GEN_214 = count >= 10'h2c & count <= 10'h33 ? 1'h0 : _GEN_189; // @[FSM.scala 268:47 FSM.scala 272:23]
  wire  _GEN_215 = count >= 10'h2c & count <= 10'h33 ? 1'h0 : _GEN_190; // @[FSM.scala 268:47 FSM.scala 272:23]
  wire  _GEN_216 = count >= 10'h2c & count <= 10'h33 ? 1'h0 : _GEN_191; // @[FSM.scala 268:47 FSM.scala 272:23]
  wire  _GEN_217 = count >= 10'h2c & count <= 10'h33 ? 1'h0 : _GEN_192; // @[FSM.scala 268:47 FSM.scala 272:23]
  wire  _GEN_218 = count >= 10'h2c & count <= 10'h33 ? 1'h0 : _GEN_193; // @[FSM.scala 268:47 FSM.scala 272:23]
  wire [9:0] _GEN_231 = count == 10'h34 ? 10'h0 : _GEN_84; // @[FSM.scala 276:27 FSM.scala 280:15]
  wire [6:0] _GEN_232 = count == 10'h34 ? 7'h0 : _GEN_85; // @[FSM.scala 276:27 FSM.scala 281:16]
  wire [2:0] _GEN_233 = count == 10'h34 ? 3'h3 : state; // @[FSM.scala 276:27 FSM.scala 282:15 FSM.scala 159:22]
  wire  _T_32 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire [9:0] _GEN_234 = count != 10'h195 ? _count_T_1 : count; // @[FSM.scala 287:28 FSM.scala 288:15 FSM.scala 161:22]
  wire [2:0] _GEN_237 = _T_3 ? 3'h2 : PEArray_ctrl_2_control; // @[FSM.scala 303:26 FSM.scala 305:33 FSM.scala 64:28]
  wire [11:0] _GEN_238 = _T_3 ? 12'h800 : PEArray_ctrl_2_mask; // @[FSM.scala 303:26 FSM.scala 306:30 FSM.scala 64:28]
  wire [11:0] _GEN_239 = _T_3 ? 12'h190 : L1_rd_addr_0; // @[FSM.scala 303:26 FSM.scala 309:25 FSM.scala 60:28]
  wire [11:0] _GEN_240 = _T_3 ? 12'h190 : L1_rd_addr_1; // @[FSM.scala 303:26 FSM.scala 309:25 FSM.scala 60:28]
  wire [11:0] _GEN_241 = _T_3 ? 12'h190 : L1_rd_addr_2; // @[FSM.scala 303:26 FSM.scala 309:25 FSM.scala 60:28]
  wire [11:0] _GEN_242 = _T_3 ? 12'h190 : L1_rd_addr_3; // @[FSM.scala 303:26 FSM.scala 309:25 FSM.scala 60:28]
  wire [11:0] _GEN_243 = _T_3 ? 12'h190 : L1_rd_addr_4; // @[FSM.scala 303:26 FSM.scala 309:25 FSM.scala 60:28]
  wire [11:0] _GEN_244 = _T_3 ? 12'h190 : L1_rd_addr_5; // @[FSM.scala 303:26 FSM.scala 309:25 FSM.scala 60:28]
  wire [11:0] _GEN_245 = _T_3 ? 12'h190 : L1_rd_addr_6; // @[FSM.scala 303:26 FSM.scala 309:25 FSM.scala 60:28]
  wire [11:0] _GEN_246 = _T_3 ? 12'h190 : L1_rd_addr_7; // @[FSM.scala 303:26 FSM.scala 309:25 FSM.scala 60:28]
  wire [11:0] _GEN_247 = _T_3 ? 12'h190 : L1_rd_addr_8; // @[FSM.scala 303:26 FSM.scala 309:25 FSM.scala 60:28]
  wire [11:0] _GEN_248 = _T_3 ? 12'h190 : L1_rd_addr_9; // @[FSM.scala 303:26 FSM.scala 309:25 FSM.scala 60:28]
  wire [11:0] _GEN_249 = _T_3 ? 12'h190 : L1_rd_addr_10; // @[FSM.scala 303:26 FSM.scala 309:25 FSM.scala 60:28]
  wire [11:0] _GEN_250 = _T_3 ? 12'h190 : L1_rd_addr_11; // @[FSM.scala 303:26 FSM.scala 309:25 FSM.scala 60:28]
  wire [11:0] _GEN_253 = _T_3 ? 12'h0 : L1_wr_addr_0; // @[FSM.scala 303:26 FSM.scala 315:25 FSM.scala 62:28]
  wire [1:0] _GEN_254 = _T_3 ? 2'h1 : BNArray_ctrl_0; // @[FSM.scala 303:26 FSM.scala 316:27 FSM.scala 65:28]
  wire  _GEN_255 = _T_3 | Relu6Array_ctrl_0; // @[FSM.scala 303:26 FSM.scala 317:30 FSM.scala 73:28]
  wire [11:0] _GEN_256 = _T_3 ? 12'h0 : L1_wr_addr_1; // @[FSM.scala 303:26 FSM.scala 315:25 FSM.scala 62:28]
  wire [1:0] _GEN_257 = _T_3 ? 2'h1 : BNArray_ctrl_1; // @[FSM.scala 303:26 FSM.scala 316:27 FSM.scala 65:28]
  wire  _GEN_258 = _T_3 | Relu6Array_ctrl_1; // @[FSM.scala 303:26 FSM.scala 317:30 FSM.scala 73:28]
  wire [11:0] _GEN_259 = _T_3 ? 12'h0 : L1_wr_addr_2; // @[FSM.scala 303:26 FSM.scala 315:25 FSM.scala 62:28]
  wire [1:0] _GEN_260 = _T_3 ? 2'h1 : BNArray_ctrl_2; // @[FSM.scala 303:26 FSM.scala 316:27 FSM.scala 65:28]
  wire  _GEN_261 = _T_3 | Relu6Array_ctrl_2; // @[FSM.scala 303:26 FSM.scala 317:30 FSM.scala 73:28]
  wire [11:0] _GEN_262 = _T_3 ? 12'h0 : L1_wr_addr_3; // @[FSM.scala 303:26 FSM.scala 315:25 FSM.scala 62:28]
  wire [1:0] _GEN_263 = _T_3 ? 2'h1 : BNArray_ctrl_3; // @[FSM.scala 303:26 FSM.scala 316:27 FSM.scala 65:28]
  wire  _GEN_264 = _T_3 | Relu6Array_ctrl_3; // @[FSM.scala 303:26 FSM.scala 317:30 FSM.scala 73:28]
  wire [11:0] _GEN_265 = _T_3 ? 12'h0 : L1_wr_addr_4; // @[FSM.scala 303:26 FSM.scala 315:25 FSM.scala 62:28]
  wire [1:0] _GEN_266 = _T_3 ? 2'h1 : BNArray_ctrl_4; // @[FSM.scala 303:26 FSM.scala 316:27 FSM.scala 65:28]
  wire  _GEN_267 = _T_3 | Relu6Array_ctrl_4; // @[FSM.scala 303:26 FSM.scala 317:30 FSM.scala 73:28]
  wire [11:0] _GEN_268 = _T_3 ? 12'h0 : L1_wr_addr_5; // @[FSM.scala 303:26 FSM.scala 315:25 FSM.scala 62:28]
  wire [1:0] _GEN_269 = _T_3 ? 2'h1 : BNArray_ctrl_5; // @[FSM.scala 303:26 FSM.scala 316:27 FSM.scala 65:28]
  wire  _GEN_270 = _T_3 | Relu6Array_ctrl_5; // @[FSM.scala 303:26 FSM.scala 317:30 FSM.scala 73:28]
  wire [11:0] _GEN_271 = _T_3 ? 12'h0 : L1_wr_addr_6; // @[FSM.scala 303:26 FSM.scala 315:25 FSM.scala 62:28]
  wire [1:0] _GEN_272 = _T_3 ? 2'h1 : BNArray_ctrl_6; // @[FSM.scala 303:26 FSM.scala 316:27 FSM.scala 65:28]
  wire  _GEN_273 = _T_3 | Relu6Array_ctrl_6; // @[FSM.scala 303:26 FSM.scala 317:30 FSM.scala 73:28]
  wire [11:0] _GEN_274 = _T_3 ? 12'h0 : L1_wr_addr_7; // @[FSM.scala 303:26 FSM.scala 315:25 FSM.scala 62:28]
  wire [1:0] _GEN_275 = _T_3 ? 2'h1 : BNArray_ctrl_7; // @[FSM.scala 303:26 FSM.scala 316:27 FSM.scala 65:28]
  wire  _GEN_276 = _T_3 | Relu6Array_ctrl_7; // @[FSM.scala 303:26 FSM.scala 317:30 FSM.scala 73:28]
  wire [11:0] _GEN_277 = _T_3 ? 12'h0 : L1_wr_addr_8; // @[FSM.scala 303:26 FSM.scala 315:25 FSM.scala 62:28]
  wire [1:0] _GEN_278 = _T_3 ? 2'h1 : BNArray_ctrl_8; // @[FSM.scala 303:26 FSM.scala 316:27 FSM.scala 65:28]
  wire  _GEN_279 = _T_3 | Relu6Array_ctrl_8; // @[FSM.scala 303:26 FSM.scala 317:30 FSM.scala 73:28]
  wire [11:0] _GEN_280 = _T_3 ? 12'h0 : L1_wr_addr_9; // @[FSM.scala 303:26 FSM.scala 315:25 FSM.scala 62:28]
  wire [1:0] _GEN_281 = _T_3 ? 2'h1 : BNArray_ctrl_9; // @[FSM.scala 303:26 FSM.scala 316:27 FSM.scala 65:28]
  wire  _GEN_282 = _T_3 | Relu6Array_ctrl_9; // @[FSM.scala 303:26 FSM.scala 317:30 FSM.scala 73:28]
  wire [11:0] _GEN_283 = _T_3 ? 12'h0 : L1_wr_addr_10; // @[FSM.scala 303:26 FSM.scala 315:25 FSM.scala 62:28]
  wire [1:0] _GEN_284 = _T_3 ? 2'h1 : BNArray_ctrl_10; // @[FSM.scala 303:26 FSM.scala 316:27 FSM.scala 65:28]
  wire  _GEN_285 = _T_3 | Relu6Array_ctrl_10; // @[FSM.scala 303:26 FSM.scala 317:30 FSM.scala 73:28]
  wire [11:0] _GEN_286 = _T_3 ? 12'h0 : L1_wr_addr_11; // @[FSM.scala 303:26 FSM.scala 315:25 FSM.scala 62:28]
  wire [1:0] _GEN_287 = _T_3 ? 2'h1 : BNArray_ctrl_11; // @[FSM.scala 303:26 FSM.scala 316:27 FSM.scala 65:28]
  wire  _GEN_288 = _T_3 | Relu6Array_ctrl_11; // @[FSM.scala 303:26 FSM.scala 317:30 FSM.scala 73:28]
  wire  _T_39 = _T_18 & count <= 10'hb; // @[FSM.scala 322:27]
  wire [2:0] _GEN_289 = _T_18 & count <= 10'hb ? 3'h2 : _GEN_237; // @[FSM.scala 322:46 FSM.scala 323:33]
  wire [11:0] _GEN_290 = _T_18 & count <= 10'hb ? {{1'd0}, PEArray_ctrl_2_mask[11:1]} : _GEN_238; // @[FSM.scala 322:46 FSM.scala 324:30]
  wire  _T_40 = count == 10'hc; // @[FSM.scala 326:18]
  wire [11:0] _GEN_291 = count == 10'hc ? 12'h0 : PEArray_ctrl_0_mask; // @[FSM.scala 326:27 FSM.scala 328:32 FSM.scala 64:28]
  wire [11:0] _GEN_292 = count == 10'hc ? 12'h0 : PEArray_ctrl_1_mask; // @[FSM.scala 326:27 FSM.scala 328:32 FSM.scala 64:28]
  wire [11:0] _GEN_293 = count == 10'hc ? 12'h0 : _GEN_290; // @[FSM.scala 326:27 FSM.scala 328:32]
  wire [11:0] _GEN_295 = 4'h1 == read_index ? L1_rd_addr_1 : L1_rd_addr_0; // @[FSM.scala 334:58 FSM.scala 334:58]
  wire [11:0] _GEN_296 = 4'h2 == read_index ? L1_rd_addr_2 : _GEN_295; // @[FSM.scala 334:58 FSM.scala 334:58]
  wire [11:0] _GEN_297 = 4'h3 == read_index ? L1_rd_addr_3 : _GEN_296; // @[FSM.scala 334:58 FSM.scala 334:58]
  wire [11:0] _GEN_298 = 4'h4 == read_index ? L1_rd_addr_4 : _GEN_297; // @[FSM.scala 334:58 FSM.scala 334:58]
  wire [11:0] _GEN_299 = 4'h5 == read_index ? L1_rd_addr_5 : _GEN_298; // @[FSM.scala 334:58 FSM.scala 334:58]
  wire [11:0] _GEN_300 = 4'h6 == read_index ? L1_rd_addr_6 : _GEN_299; // @[FSM.scala 334:58 FSM.scala 334:58]
  wire [11:0] _GEN_301 = 4'h7 == read_index ? L1_rd_addr_7 : _GEN_300; // @[FSM.scala 334:58 FSM.scala 334:58]
  wire [11:0] _GEN_302 = 4'h8 == read_index ? L1_rd_addr_8 : _GEN_301; // @[FSM.scala 334:58 FSM.scala 334:58]
  wire [11:0] _GEN_303 = 4'h9 == read_index ? L1_rd_addr_9 : _GEN_302; // @[FSM.scala 334:58 FSM.scala 334:58]
  wire [11:0] _GEN_304 = 4'ha == read_index ? L1_rd_addr_10 : _GEN_303; // @[FSM.scala 334:58 FSM.scala 334:58]
  wire [11:0] _GEN_305 = 4'hb == read_index ? L1_rd_addr_11 : _GEN_304; // @[FSM.scala 334:58 FSM.scala 334:58]
  wire [11:0] _L1_rd_addr_T_1 = _GEN_305 + 12'h1; // @[FSM.scala 334:58]
  wire [11:0] _GEN_306 = 4'h0 == read_index ? _L1_rd_addr_T_1 : _GEN_239; // @[FSM.scala 334:32 FSM.scala 334:32]
  wire [11:0] _GEN_307 = 4'h1 == read_index ? _L1_rd_addr_T_1 : _GEN_240; // @[FSM.scala 334:32 FSM.scala 334:32]
  wire [11:0] _GEN_308 = 4'h2 == read_index ? _L1_rd_addr_T_1 : _GEN_241; // @[FSM.scala 334:32 FSM.scala 334:32]
  wire [11:0] _GEN_309 = 4'h3 == read_index ? _L1_rd_addr_T_1 : _GEN_242; // @[FSM.scala 334:32 FSM.scala 334:32]
  wire [11:0] _GEN_310 = 4'h4 == read_index ? _L1_rd_addr_T_1 : _GEN_243; // @[FSM.scala 334:32 FSM.scala 334:32]
  wire [11:0] _GEN_311 = 4'h5 == read_index ? _L1_rd_addr_T_1 : _GEN_244; // @[FSM.scala 334:32 FSM.scala 334:32]
  wire [11:0] _GEN_312 = 4'h6 == read_index ? _L1_rd_addr_T_1 : _GEN_245; // @[FSM.scala 334:32 FSM.scala 334:32]
  wire [11:0] _GEN_313 = 4'h7 == read_index ? _L1_rd_addr_T_1 : _GEN_246; // @[FSM.scala 334:32 FSM.scala 334:32]
  wire [11:0] _GEN_314 = 4'h8 == read_index ? _L1_rd_addr_T_1 : _GEN_247; // @[FSM.scala 334:32 FSM.scala 334:32]
  wire [11:0] _GEN_315 = 4'h9 == read_index ? _L1_rd_addr_T_1 : _GEN_248; // @[FSM.scala 334:32 FSM.scala 334:32]
  wire [11:0] _GEN_316 = 4'ha == read_index ? _L1_rd_addr_T_1 : _GEN_249; // @[FSM.scala 334:32 FSM.scala 334:32]
  wire [11:0] _GEN_317 = 4'hb == read_index ? _L1_rd_addr_T_1 : _GEN_250; // @[FSM.scala 334:32 FSM.scala 334:32]
  wire [3:0] _read_index_T_1 = read_index + 4'h1; // @[FSM.scala 336:36]
  wire [3:0] _PE_rd_data_mux_T_1 = PE_rd_data_mux + 4'h1; // @[FSM.scala 337:44]
  wire [3:0] _GEN_318 = count1 == 7'h7 ? _read_index_T_1 : read_index; // @[FSM.scala 335:52 FSM.scala 336:22 FSM.scala 165:27]
  wire [3:0] _GEN_319 = count1 == 7'h7 ? _PE_rd_data_mux_T_1 : _GEN_105; // @[FSM.scala 335:52 FSM.scala 337:26]
  wire [11:0] _GEN_321 = _T_18 & count <= 10'h187 ? _GEN_306 : _GEN_239; // @[FSM.scala 333:43]
  wire [11:0] _GEN_322 = _T_18 & count <= 10'h187 ? _GEN_307 : _GEN_240; // @[FSM.scala 333:43]
  wire [11:0] _GEN_323 = _T_18 & count <= 10'h187 ? _GEN_308 : _GEN_241; // @[FSM.scala 333:43]
  wire [11:0] _GEN_324 = _T_18 & count <= 10'h187 ? _GEN_309 : _GEN_242; // @[FSM.scala 333:43]
  wire [11:0] _GEN_325 = _T_18 & count <= 10'h187 ? _GEN_310 : _GEN_243; // @[FSM.scala 333:43]
  wire [11:0] _GEN_326 = _T_18 & count <= 10'h187 ? _GEN_311 : _GEN_244; // @[FSM.scala 333:43]
  wire [11:0] _GEN_327 = _T_18 & count <= 10'h187 ? _GEN_312 : _GEN_245; // @[FSM.scala 333:43]
  wire [11:0] _GEN_328 = _T_18 & count <= 10'h187 ? _GEN_313 : _GEN_246; // @[FSM.scala 333:43]
  wire [11:0] _GEN_329 = _T_18 & count <= 10'h187 ? _GEN_314 : _GEN_247; // @[FSM.scala 333:43]
  wire [11:0] _GEN_330 = _T_18 & count <= 10'h187 ? _GEN_315 : _GEN_248; // @[FSM.scala 333:43]
  wire [11:0] _GEN_331 = _T_18 & count <= 10'h187 ? _GEN_316 : _GEN_249; // @[FSM.scala 333:43]
  wire [11:0] _GEN_332 = _T_18 & count <= 10'h187 ? _GEN_317 : _GEN_250; // @[FSM.scala 333:43]
  wire [3:0] _GEN_333 = _T_18 & count <= 10'h187 ? _GEN_318 : read_index; // @[FSM.scala 333:43 FSM.scala 165:27]
  wire [3:0] _GEN_334 = _T_18 & count <= 10'h187 ? _GEN_319 : _GEN_105; // @[FSM.scala 333:43]
  wire  _T_48 = count == 10'h2; // @[FSM.scala 345:18]
  wire  _GEN_335 = count == 10'h2 | L1_wrEna_0; // @[FSM.scala 345:26 FSM.scala 347:23 FSM.scala 63:28]
  wire [11:0] _GEN_336 = count == 10'h2 ? _L1_wr_addr_0_T_1 : _GEN_253; // @[FSM.scala 345:26 FSM.scala 348:25]
  wire  _T_49 = count == 10'h3; // @[FSM.scala 351:18]
  wire  _GEN_337 = count == 10'h3 | _GEN_335; // @[FSM.scala 351:26 FSM.scala 353:23]
  wire [11:0] _GEN_338 = count == 10'h3 ? _L1_wr_addr_0_T_1 : _GEN_336; // @[FSM.scala 351:26 FSM.scala 354:25]
  wire  _GEN_339 = count == 10'h3 | L1_wrEna_1; // @[FSM.scala 351:26 FSM.scala 353:23 FSM.scala 63:28]
  wire [11:0] _GEN_340 = count == 10'h3 ? _L1_wr_addr_1_T_1 : _GEN_256; // @[FSM.scala 351:26 FSM.scala 354:25]
  wire  _GEN_341 = _T_21 | _GEN_337; // @[FSM.scala 357:26 FSM.scala 359:23]
  wire [11:0] _GEN_342 = _T_21 ? _L1_wr_addr_0_T_1 : _GEN_338; // @[FSM.scala 357:26 FSM.scala 360:25]
  wire  _GEN_343 = _T_21 | _GEN_339; // @[FSM.scala 357:26 FSM.scala 359:23]
  wire [11:0] _GEN_344 = _T_21 ? _L1_wr_addr_1_T_1 : _GEN_340; // @[FSM.scala 357:26 FSM.scala 360:25]
  wire [11:0] _GEN_346 = _T_21 ? _L1_wr_addr_2_T_1 : _GEN_259; // @[FSM.scala 357:26 FSM.scala 360:25]
  wire  _T_51 = count == 10'h5; // @[FSM.scala 363:18]
  wire  _GEN_347 = count == 10'h5 | _GEN_341; // @[FSM.scala 363:26 FSM.scala 365:23]
  wire [11:0] _GEN_348 = count == 10'h5 ? _L1_wr_addr_0_T_1 : _GEN_342; // @[FSM.scala 363:26 FSM.scala 366:25]
  wire  _GEN_349 = count == 10'h5 | _GEN_343; // @[FSM.scala 363:26 FSM.scala 365:23]
  wire [11:0] _GEN_350 = count == 10'h5 ? _L1_wr_addr_1_T_1 : _GEN_344; // @[FSM.scala 363:26 FSM.scala 366:25]
  wire  _GEN_351 = count == 10'h5 | _GEN_129; // @[FSM.scala 363:26 FSM.scala 365:23]
  wire [11:0] _GEN_352 = count == 10'h5 ? _L1_wr_addr_2_T_1 : _GEN_346; // @[FSM.scala 363:26 FSM.scala 366:25]
  wire  _GEN_353 = count == 10'h5 | L1_wrEna_3; // @[FSM.scala 363:26 FSM.scala 365:23 FSM.scala 63:28]
  wire [11:0] _GEN_354 = count == 10'h5 ? _L1_wr_addr_3_T_1 : _GEN_262; // @[FSM.scala 363:26 FSM.scala 366:25]
  wire  _T_52 = count == 10'h6; // @[FSM.scala 369:18]
  wire  _GEN_355 = count == 10'h6 | _GEN_347; // @[FSM.scala 369:26 FSM.scala 371:23]
  wire [11:0] _GEN_356 = count == 10'h6 ? _L1_wr_addr_0_T_1 : _GEN_348; // @[FSM.scala 369:26 FSM.scala 372:25]
  wire  _GEN_357 = count == 10'h6 | _GEN_349; // @[FSM.scala 369:26 FSM.scala 371:23]
  wire [11:0] _GEN_358 = count == 10'h6 ? _L1_wr_addr_1_T_1 : _GEN_350; // @[FSM.scala 369:26 FSM.scala 372:25]
  wire  _GEN_359 = count == 10'h6 | _GEN_351; // @[FSM.scala 369:26 FSM.scala 371:23]
  wire [11:0] _GEN_360 = count == 10'h6 ? _L1_wr_addr_2_T_1 : _GEN_352; // @[FSM.scala 369:26 FSM.scala 372:25]
  wire  _GEN_361 = count == 10'h6 | _GEN_353; // @[FSM.scala 369:26 FSM.scala 371:23]
  wire [11:0] _GEN_362 = count == 10'h6 ? _L1_wr_addr_3_T_1 : _GEN_354; // @[FSM.scala 369:26 FSM.scala 372:25]
  wire  _GEN_363 = count == 10'h6 | L1_wrEna_4; // @[FSM.scala 369:26 FSM.scala 371:23 FSM.scala 63:28]
  wire [11:0] _GEN_364 = count == 10'h6 ? _L1_wr_addr_4_T_1 : _GEN_265; // @[FSM.scala 369:26 FSM.scala 372:25]
  wire  _T_53 = count == 10'h7; // @[FSM.scala 375:18]
  wire  _GEN_365 = count == 10'h7 | _GEN_355; // @[FSM.scala 375:26 FSM.scala 377:23]
  wire [11:0] _GEN_366 = count == 10'h7 ? _L1_wr_addr_0_T_1 : _GEN_356; // @[FSM.scala 375:26 FSM.scala 378:25]
  wire  _GEN_367 = count == 10'h7 | _GEN_357; // @[FSM.scala 375:26 FSM.scala 377:23]
  wire [11:0] _GEN_368 = count == 10'h7 ? _L1_wr_addr_1_T_1 : _GEN_358; // @[FSM.scala 375:26 FSM.scala 378:25]
  wire  _GEN_369 = count == 10'h7 | _GEN_359; // @[FSM.scala 375:26 FSM.scala 377:23]
  wire [11:0] _GEN_370 = count == 10'h7 ? _L1_wr_addr_2_T_1 : _GEN_360; // @[FSM.scala 375:26 FSM.scala 378:25]
  wire  _GEN_371 = count == 10'h7 | _GEN_361; // @[FSM.scala 375:26 FSM.scala 377:23]
  wire [11:0] _GEN_372 = count == 10'h7 ? _L1_wr_addr_3_T_1 : _GEN_362; // @[FSM.scala 375:26 FSM.scala 378:25]
  wire  _GEN_373 = count == 10'h7 | _GEN_363; // @[FSM.scala 375:26 FSM.scala 377:23]
  wire [11:0] _GEN_374 = count == 10'h7 ? _L1_wr_addr_4_T_1 : _GEN_364; // @[FSM.scala 375:26 FSM.scala 378:25]
  wire  _GEN_375 = count == 10'h7 | L1_wrEna_5; // @[FSM.scala 375:26 FSM.scala 377:23 FSM.scala 63:28]
  wire [11:0] _GEN_376 = count == 10'h7 ? _L1_wr_addr_5_T_1 : _GEN_268; // @[FSM.scala 375:26 FSM.scala 378:25]
  wire  _T_54 = count == 10'h8; // @[FSM.scala 381:18]
  wire  _GEN_377 = count == 10'h8 | _GEN_365; // @[FSM.scala 381:26 FSM.scala 383:23]
  wire [11:0] _GEN_378 = count == 10'h8 ? _L1_wr_addr_0_T_1 : _GEN_366; // @[FSM.scala 381:26 FSM.scala 384:25]
  wire  _GEN_379 = count == 10'h8 | _GEN_367; // @[FSM.scala 381:26 FSM.scala 383:23]
  wire [11:0] _GEN_380 = count == 10'h8 ? _L1_wr_addr_1_T_1 : _GEN_368; // @[FSM.scala 381:26 FSM.scala 384:25]
  wire  _GEN_381 = count == 10'h8 | _GEN_369; // @[FSM.scala 381:26 FSM.scala 383:23]
  wire [11:0] _GEN_382 = count == 10'h8 ? _L1_wr_addr_2_T_1 : _GEN_370; // @[FSM.scala 381:26 FSM.scala 384:25]
  wire  _GEN_383 = count == 10'h8 | _GEN_371; // @[FSM.scala 381:26 FSM.scala 383:23]
  wire [11:0] _GEN_384 = count == 10'h8 ? _L1_wr_addr_3_T_1 : _GEN_372; // @[FSM.scala 381:26 FSM.scala 384:25]
  wire  _GEN_385 = count == 10'h8 | _GEN_373; // @[FSM.scala 381:26 FSM.scala 383:23]
  wire [11:0] _GEN_386 = count == 10'h8 ? _L1_wr_addr_4_T_1 : _GEN_374; // @[FSM.scala 381:26 FSM.scala 384:25]
  wire  _GEN_387 = count == 10'h8 | _GEN_375; // @[FSM.scala 381:26 FSM.scala 383:23]
  wire [11:0] _GEN_388 = count == 10'h8 ? _L1_wr_addr_5_T_1 : _GEN_376; // @[FSM.scala 381:26 FSM.scala 384:25]
  wire  _GEN_389 = count == 10'h8 | L1_wrEna_6; // @[FSM.scala 381:26 FSM.scala 383:23 FSM.scala 63:28]
  wire [11:0] _GEN_390 = count == 10'h8 ? _L1_wr_addr_6_T_1 : _GEN_271; // @[FSM.scala 381:26 FSM.scala 384:25]
  wire  _T_55 = count == 10'h9; // @[FSM.scala 387:18]
  wire  _GEN_391 = count == 10'h9 | _GEN_377; // @[FSM.scala 387:26 FSM.scala 389:23]
  wire [11:0] _GEN_392 = count == 10'h9 ? _L1_wr_addr_0_T_1 : _GEN_378; // @[FSM.scala 387:26 FSM.scala 390:25]
  wire  _GEN_393 = count == 10'h9 | _GEN_379; // @[FSM.scala 387:26 FSM.scala 389:23]
  wire [11:0] _GEN_394 = count == 10'h9 ? _L1_wr_addr_1_T_1 : _GEN_380; // @[FSM.scala 387:26 FSM.scala 390:25]
  wire  _GEN_395 = count == 10'h9 | _GEN_381; // @[FSM.scala 387:26 FSM.scala 389:23]
  wire [11:0] _GEN_396 = count == 10'h9 ? _L1_wr_addr_2_T_1 : _GEN_382; // @[FSM.scala 387:26 FSM.scala 390:25]
  wire  _GEN_397 = count == 10'h9 | _GEN_383; // @[FSM.scala 387:26 FSM.scala 389:23]
  wire [11:0] _GEN_398 = count == 10'h9 ? _L1_wr_addr_3_T_1 : _GEN_384; // @[FSM.scala 387:26 FSM.scala 390:25]
  wire  _GEN_399 = count == 10'h9 | _GEN_385; // @[FSM.scala 387:26 FSM.scala 389:23]
  wire [11:0] _GEN_400 = count == 10'h9 ? _L1_wr_addr_4_T_1 : _GEN_386; // @[FSM.scala 387:26 FSM.scala 390:25]
  wire  _GEN_401 = count == 10'h9 | _GEN_387; // @[FSM.scala 387:26 FSM.scala 389:23]
  wire [11:0] _GEN_402 = count == 10'h9 ? _L1_wr_addr_5_T_1 : _GEN_388; // @[FSM.scala 387:26 FSM.scala 390:25]
  wire  _GEN_403 = count == 10'h9 | _GEN_389; // @[FSM.scala 387:26 FSM.scala 389:23]
  wire [11:0] _GEN_404 = count == 10'h9 ? _L1_wr_addr_6_T_1 : _GEN_390; // @[FSM.scala 387:26 FSM.scala 390:25]
  wire  _GEN_405 = count == 10'h9 | L1_wrEna_7; // @[FSM.scala 387:26 FSM.scala 389:23 FSM.scala 63:28]
  wire [11:0] _GEN_406 = count == 10'h9 ? _L1_wr_addr_7_T_1 : _GEN_274; // @[FSM.scala 387:26 FSM.scala 390:25]
  wire  _T_56 = count == 10'ha; // @[FSM.scala 393:18]
  wire  _GEN_407 = count == 10'ha | _GEN_391; // @[FSM.scala 393:27 FSM.scala 395:23]
  wire [11:0] _GEN_408 = count == 10'ha ? _L1_wr_addr_0_T_1 : _GEN_392; // @[FSM.scala 393:27 FSM.scala 396:25]
  wire  _GEN_409 = count == 10'ha | _GEN_393; // @[FSM.scala 393:27 FSM.scala 395:23]
  wire [11:0] _GEN_410 = count == 10'ha ? _L1_wr_addr_1_T_1 : _GEN_394; // @[FSM.scala 393:27 FSM.scala 396:25]
  wire  _GEN_411 = count == 10'ha | _GEN_395; // @[FSM.scala 393:27 FSM.scala 395:23]
  wire [11:0] _GEN_412 = count == 10'ha ? _L1_wr_addr_2_T_1 : _GEN_396; // @[FSM.scala 393:27 FSM.scala 396:25]
  wire  _GEN_413 = count == 10'ha | _GEN_397; // @[FSM.scala 393:27 FSM.scala 395:23]
  wire [11:0] _GEN_414 = count == 10'ha ? _L1_wr_addr_3_T_1 : _GEN_398; // @[FSM.scala 393:27 FSM.scala 396:25]
  wire  _GEN_415 = count == 10'ha | _GEN_399; // @[FSM.scala 393:27 FSM.scala 395:23]
  wire [11:0] _GEN_416 = count == 10'ha ? _L1_wr_addr_4_T_1 : _GEN_400; // @[FSM.scala 393:27 FSM.scala 396:25]
  wire  _GEN_417 = count == 10'ha | _GEN_401; // @[FSM.scala 393:27 FSM.scala 395:23]
  wire [11:0] _GEN_418 = count == 10'ha ? _L1_wr_addr_5_T_1 : _GEN_402; // @[FSM.scala 393:27 FSM.scala 396:25]
  wire  _GEN_419 = count == 10'ha | _GEN_403; // @[FSM.scala 393:27 FSM.scala 395:23]
  wire [11:0] _GEN_420 = count == 10'ha ? _L1_wr_addr_6_T_1 : _GEN_404; // @[FSM.scala 393:27 FSM.scala 396:25]
  wire  _GEN_421 = count == 10'ha | _GEN_405; // @[FSM.scala 393:27 FSM.scala 395:23]
  wire [11:0] _GEN_422 = count == 10'ha ? _L1_wr_addr_7_T_1 : _GEN_406; // @[FSM.scala 393:27 FSM.scala 396:25]
  wire  _GEN_423 = count == 10'ha | L1_wrEna_8; // @[FSM.scala 393:27 FSM.scala 395:23 FSM.scala 63:28]
  wire [11:0] _GEN_424 = count == 10'ha ? _L1_wr_addr_8_T_1 : _GEN_277; // @[FSM.scala 393:27 FSM.scala 396:25]
  wire  _T_57 = count == 10'hb; // @[FSM.scala 399:18]
  wire  _GEN_425 = count == 10'hb | _GEN_407; // @[FSM.scala 399:27 FSM.scala 401:23]
  wire [11:0] _GEN_426 = count == 10'hb ? _L1_wr_addr_0_T_1 : _GEN_408; // @[FSM.scala 399:27 FSM.scala 402:25]
  wire  _GEN_427 = count == 10'hb | _GEN_409; // @[FSM.scala 399:27 FSM.scala 401:23]
  wire [11:0] _GEN_428 = count == 10'hb ? _L1_wr_addr_1_T_1 : _GEN_410; // @[FSM.scala 399:27 FSM.scala 402:25]
  wire  _GEN_429 = count == 10'hb | _GEN_411; // @[FSM.scala 399:27 FSM.scala 401:23]
  wire [11:0] _GEN_430 = count == 10'hb ? _L1_wr_addr_2_T_1 : _GEN_412; // @[FSM.scala 399:27 FSM.scala 402:25]
  wire  _GEN_431 = count == 10'hb | _GEN_413; // @[FSM.scala 399:27 FSM.scala 401:23]
  wire [11:0] _GEN_432 = count == 10'hb ? _L1_wr_addr_3_T_1 : _GEN_414; // @[FSM.scala 399:27 FSM.scala 402:25]
  wire  _GEN_433 = count == 10'hb | _GEN_415; // @[FSM.scala 399:27 FSM.scala 401:23]
  wire [11:0] _GEN_434 = count == 10'hb ? _L1_wr_addr_4_T_1 : _GEN_416; // @[FSM.scala 399:27 FSM.scala 402:25]
  wire  _GEN_435 = count == 10'hb | _GEN_417; // @[FSM.scala 399:27 FSM.scala 401:23]
  wire [11:0] _GEN_436 = count == 10'hb ? _L1_wr_addr_5_T_1 : _GEN_418; // @[FSM.scala 399:27 FSM.scala 402:25]
  wire  _GEN_437 = count == 10'hb | _GEN_419; // @[FSM.scala 399:27 FSM.scala 401:23]
  wire [11:0] _GEN_438 = count == 10'hb ? _L1_wr_addr_6_T_1 : _GEN_420; // @[FSM.scala 399:27 FSM.scala 402:25]
  wire  _GEN_439 = count == 10'hb | _GEN_421; // @[FSM.scala 399:27 FSM.scala 401:23]
  wire [11:0] _GEN_440 = count == 10'hb ? _L1_wr_addr_7_T_1 : _GEN_422; // @[FSM.scala 399:27 FSM.scala 402:25]
  wire  _GEN_441 = count == 10'hb | _GEN_423; // @[FSM.scala 399:27 FSM.scala 401:23]
  wire [11:0] _GEN_442 = count == 10'hb ? _L1_wr_addr_8_T_1 : _GEN_424; // @[FSM.scala 399:27 FSM.scala 402:25]
  wire  _GEN_443 = count == 10'hb | L1_wrEna_9; // @[FSM.scala 399:27 FSM.scala 401:23 FSM.scala 63:28]
  wire [11:0] _GEN_444 = count == 10'hb ? _L1_wr_addr_9_T_1 : _GEN_280; // @[FSM.scala 399:27 FSM.scala 402:25]
  wire  _GEN_445 = _T_40 | _GEN_425; // @[FSM.scala 405:27 FSM.scala 407:23]
  wire [11:0] _GEN_446 = _T_40 ? _L1_wr_addr_0_T_1 : _GEN_426; // @[FSM.scala 405:27 FSM.scala 408:25]
  wire  _GEN_447 = _T_40 | _GEN_427; // @[FSM.scala 405:27 FSM.scala 407:23]
  wire [11:0] _GEN_448 = _T_40 ? _L1_wr_addr_1_T_1 : _GEN_428; // @[FSM.scala 405:27 FSM.scala 408:25]
  wire  _GEN_449 = _T_40 | _GEN_429; // @[FSM.scala 405:27 FSM.scala 407:23]
  wire [11:0] _GEN_450 = _T_40 ? _L1_wr_addr_2_T_1 : _GEN_430; // @[FSM.scala 405:27 FSM.scala 408:25]
  wire  _GEN_451 = _T_40 | _GEN_431; // @[FSM.scala 405:27 FSM.scala 407:23]
  wire [11:0] _GEN_452 = _T_40 ? _L1_wr_addr_3_T_1 : _GEN_432; // @[FSM.scala 405:27 FSM.scala 408:25]
  wire  _GEN_453 = _T_40 | _GEN_433; // @[FSM.scala 405:27 FSM.scala 407:23]
  wire [11:0] _GEN_454 = _T_40 ? _L1_wr_addr_4_T_1 : _GEN_434; // @[FSM.scala 405:27 FSM.scala 408:25]
  wire  _GEN_455 = _T_40 | _GEN_435; // @[FSM.scala 405:27 FSM.scala 407:23]
  wire [11:0] _GEN_456 = _T_40 ? _L1_wr_addr_5_T_1 : _GEN_436; // @[FSM.scala 405:27 FSM.scala 408:25]
  wire  _GEN_457 = _T_40 | _GEN_437; // @[FSM.scala 405:27 FSM.scala 407:23]
  wire [11:0] _GEN_458 = _T_40 ? _L1_wr_addr_6_T_1 : _GEN_438; // @[FSM.scala 405:27 FSM.scala 408:25]
  wire  _GEN_459 = _T_40 | _GEN_439; // @[FSM.scala 405:27 FSM.scala 407:23]
  wire [11:0] _GEN_460 = _T_40 ? _L1_wr_addr_7_T_1 : _GEN_440; // @[FSM.scala 405:27 FSM.scala 408:25]
  wire  _GEN_461 = _T_40 | _GEN_441; // @[FSM.scala 405:27 FSM.scala 407:23]
  wire [11:0] _GEN_462 = _T_40 ? _L1_wr_addr_8_T_1 : _GEN_442; // @[FSM.scala 405:27 FSM.scala 408:25]
  wire  _GEN_463 = _T_40 | _GEN_443; // @[FSM.scala 405:27 FSM.scala 407:23]
  wire [11:0] _GEN_464 = _T_40 ? _L1_wr_addr_9_T_1 : _GEN_444; // @[FSM.scala 405:27 FSM.scala 408:25]
  wire  _GEN_465 = _T_40 | L1_wrEna_10; // @[FSM.scala 405:27 FSM.scala 407:23 FSM.scala 63:28]
  wire [11:0] _GEN_466 = _T_40 ? _L1_wr_addr_10_T_1 : _GEN_283; // @[FSM.scala 405:27 FSM.scala 408:25]
  wire  _GEN_467 = count >= 10'hd & count <= 10'h189 | _GEN_445; // @[FSM.scala 411:48 FSM.scala 413:23]
  wire [11:0] _GEN_468 = count >= 10'hd & count <= 10'h189 ? _L1_wr_addr_0_T_1 : _GEN_446; // @[FSM.scala 411:48 FSM.scala 414:25]
  wire  _GEN_469 = count >= 10'hd & count <= 10'h189 | _GEN_447; // @[FSM.scala 411:48 FSM.scala 413:23]
  wire [11:0] _GEN_470 = count >= 10'hd & count <= 10'h189 ? _L1_wr_addr_1_T_1 : _GEN_448; // @[FSM.scala 411:48 FSM.scala 414:25]
  wire  _GEN_471 = count >= 10'hd & count <= 10'h189 | _GEN_449; // @[FSM.scala 411:48 FSM.scala 413:23]
  wire [11:0] _GEN_472 = count >= 10'hd & count <= 10'h189 ? _L1_wr_addr_2_T_1 : _GEN_450; // @[FSM.scala 411:48 FSM.scala 414:25]
  wire  _GEN_473 = count >= 10'hd & count <= 10'h189 | _GEN_451; // @[FSM.scala 411:48 FSM.scala 413:23]
  wire [11:0] _GEN_474 = count >= 10'hd & count <= 10'h189 ? _L1_wr_addr_3_T_1 : _GEN_452; // @[FSM.scala 411:48 FSM.scala 414:25]
  wire  _GEN_475 = count >= 10'hd & count <= 10'h189 | _GEN_453; // @[FSM.scala 411:48 FSM.scala 413:23]
  wire [11:0] _GEN_476 = count >= 10'hd & count <= 10'h189 ? _L1_wr_addr_4_T_1 : _GEN_454; // @[FSM.scala 411:48 FSM.scala 414:25]
  wire  _GEN_477 = count >= 10'hd & count <= 10'h189 | _GEN_455; // @[FSM.scala 411:48 FSM.scala 413:23]
  wire [11:0] _GEN_478 = count >= 10'hd & count <= 10'h189 ? _L1_wr_addr_5_T_1 : _GEN_456; // @[FSM.scala 411:48 FSM.scala 414:25]
  wire  _GEN_479 = count >= 10'hd & count <= 10'h189 | _GEN_457; // @[FSM.scala 411:48 FSM.scala 413:23]
  wire [11:0] _GEN_480 = count >= 10'hd & count <= 10'h189 ? _L1_wr_addr_6_T_1 : _GEN_458; // @[FSM.scala 411:48 FSM.scala 414:25]
  wire  _GEN_481 = count >= 10'hd & count <= 10'h189 | _GEN_459; // @[FSM.scala 411:48 FSM.scala 413:23]
  wire [11:0] _GEN_482 = count >= 10'hd & count <= 10'h189 ? _L1_wr_addr_7_T_1 : _GEN_460; // @[FSM.scala 411:48 FSM.scala 414:25]
  wire  _GEN_483 = count >= 10'hd & count <= 10'h189 | _GEN_461; // @[FSM.scala 411:48 FSM.scala 413:23]
  wire [11:0] _GEN_484 = count >= 10'hd & count <= 10'h189 ? _L1_wr_addr_8_T_1 : _GEN_462; // @[FSM.scala 411:48 FSM.scala 414:25]
  wire  _GEN_485 = count >= 10'hd & count <= 10'h189 | _GEN_463; // @[FSM.scala 411:48 FSM.scala 413:23]
  wire [11:0] _GEN_486 = count >= 10'hd & count <= 10'h189 ? _L1_wr_addr_9_T_1 : _GEN_464; // @[FSM.scala 411:48 FSM.scala 414:25]
  wire  _GEN_487 = count >= 10'hd & count <= 10'h189 | _GEN_465; // @[FSM.scala 411:48 FSM.scala 413:23]
  wire [11:0] _GEN_488 = count >= 10'hd & count <= 10'h189 ? _L1_wr_addr_10_T_1 : _GEN_466; // @[FSM.scala 411:48 FSM.scala 414:25]
  wire  _GEN_489 = count >= 10'hd & count <= 10'h189 | L1_wrEna_11; // @[FSM.scala 411:48 FSM.scala 413:23 FSM.scala 63:28]
  wire [11:0] _GEN_490 = count >= 10'hd & count <= 10'h189 ? _L1_wr_addr_11_T_1 : _GEN_286; // @[FSM.scala 411:48 FSM.scala 414:25]
  wire  _T_65 = count == 10'h18a; // @[FSM.scala 417:18]
  wire  _GEN_491 = count == 10'h18a | _GEN_469; // @[FSM.scala 417:28 FSM.scala 419:23]
  wire [11:0] _GEN_492 = count == 10'h18a ? _L1_wr_addr_1_T_1 : _GEN_470; // @[FSM.scala 417:28 FSM.scala 420:25]
  wire  _GEN_493 = count == 10'h18a | _GEN_471; // @[FSM.scala 417:28 FSM.scala 419:23]
  wire [11:0] _GEN_494 = count == 10'h18a ? _L1_wr_addr_2_T_1 : _GEN_472; // @[FSM.scala 417:28 FSM.scala 420:25]
  wire  _GEN_495 = count == 10'h18a | _GEN_473; // @[FSM.scala 417:28 FSM.scala 419:23]
  wire [11:0] _GEN_496 = count == 10'h18a ? _L1_wr_addr_3_T_1 : _GEN_474; // @[FSM.scala 417:28 FSM.scala 420:25]
  wire  _GEN_497 = count == 10'h18a | _GEN_475; // @[FSM.scala 417:28 FSM.scala 419:23]
  wire [11:0] _GEN_498 = count == 10'h18a ? _L1_wr_addr_4_T_1 : _GEN_476; // @[FSM.scala 417:28 FSM.scala 420:25]
  wire  _GEN_499 = count == 10'h18a | _GEN_477; // @[FSM.scala 417:28 FSM.scala 419:23]
  wire [11:0] _GEN_500 = count == 10'h18a ? _L1_wr_addr_5_T_1 : _GEN_478; // @[FSM.scala 417:28 FSM.scala 420:25]
  wire  _GEN_501 = count == 10'h18a | _GEN_479; // @[FSM.scala 417:28 FSM.scala 419:23]
  wire [11:0] _GEN_502 = count == 10'h18a ? _L1_wr_addr_6_T_1 : _GEN_480; // @[FSM.scala 417:28 FSM.scala 420:25]
  wire  _GEN_503 = count == 10'h18a | _GEN_481; // @[FSM.scala 417:28 FSM.scala 419:23]
  wire [11:0] _GEN_504 = count == 10'h18a ? _L1_wr_addr_7_T_1 : _GEN_482; // @[FSM.scala 417:28 FSM.scala 420:25]
  wire  _GEN_505 = count == 10'h18a | _GEN_483; // @[FSM.scala 417:28 FSM.scala 419:23]
  wire [11:0] _GEN_506 = count == 10'h18a ? _L1_wr_addr_8_T_1 : _GEN_484; // @[FSM.scala 417:28 FSM.scala 420:25]
  wire  _GEN_507 = count == 10'h18a | _GEN_485; // @[FSM.scala 417:28 FSM.scala 419:23]
  wire [11:0] _GEN_508 = count == 10'h18a ? _L1_wr_addr_9_T_1 : _GEN_486; // @[FSM.scala 417:28 FSM.scala 420:25]
  wire  _GEN_509 = count == 10'h18a | _GEN_487; // @[FSM.scala 417:28 FSM.scala 419:23]
  wire [11:0] _GEN_510 = count == 10'h18a ? _L1_wr_addr_10_T_1 : _GEN_488; // @[FSM.scala 417:28 FSM.scala 420:25]
  wire  _GEN_511 = count == 10'h18a | _GEN_489; // @[FSM.scala 417:28 FSM.scala 419:23]
  wire [11:0] _GEN_512 = count == 10'h18a ? _L1_wr_addr_11_T_1 : _GEN_490; // @[FSM.scala 417:28 FSM.scala 420:25]
  wire  _GEN_513 = count == 10'h18b | _GEN_493; // @[FSM.scala 423:28 FSM.scala 425:23]
  wire [11:0] _GEN_514 = count == 10'h18b ? _L1_wr_addr_2_T_1 : _GEN_494; // @[FSM.scala 423:28 FSM.scala 426:25]
  wire  _GEN_515 = count == 10'h18b | _GEN_495; // @[FSM.scala 423:28 FSM.scala 425:23]
  wire [11:0] _GEN_516 = count == 10'h18b ? _L1_wr_addr_3_T_1 : _GEN_496; // @[FSM.scala 423:28 FSM.scala 426:25]
  wire  _GEN_517 = count == 10'h18b | _GEN_497; // @[FSM.scala 423:28 FSM.scala 425:23]
  wire [11:0] _GEN_518 = count == 10'h18b ? _L1_wr_addr_4_T_1 : _GEN_498; // @[FSM.scala 423:28 FSM.scala 426:25]
  wire  _GEN_519 = count == 10'h18b | _GEN_499; // @[FSM.scala 423:28 FSM.scala 425:23]
  wire [11:0] _GEN_520 = count == 10'h18b ? _L1_wr_addr_5_T_1 : _GEN_500; // @[FSM.scala 423:28 FSM.scala 426:25]
  wire  _GEN_521 = count == 10'h18b | _GEN_501; // @[FSM.scala 423:28 FSM.scala 425:23]
  wire [11:0] _GEN_522 = count == 10'h18b ? _L1_wr_addr_6_T_1 : _GEN_502; // @[FSM.scala 423:28 FSM.scala 426:25]
  wire  _GEN_523 = count == 10'h18b | _GEN_503; // @[FSM.scala 423:28 FSM.scala 425:23]
  wire [11:0] _GEN_524 = count == 10'h18b ? _L1_wr_addr_7_T_1 : _GEN_504; // @[FSM.scala 423:28 FSM.scala 426:25]
  wire  _GEN_525 = count == 10'h18b | _GEN_505; // @[FSM.scala 423:28 FSM.scala 425:23]
  wire [11:0] _GEN_526 = count == 10'h18b ? _L1_wr_addr_8_T_1 : _GEN_506; // @[FSM.scala 423:28 FSM.scala 426:25]
  wire  _GEN_527 = count == 10'h18b | _GEN_507; // @[FSM.scala 423:28 FSM.scala 425:23]
  wire [11:0] _GEN_528 = count == 10'h18b ? _L1_wr_addr_9_T_1 : _GEN_508; // @[FSM.scala 423:28 FSM.scala 426:25]
  wire  _GEN_529 = count == 10'h18b | _GEN_509; // @[FSM.scala 423:28 FSM.scala 425:23]
  wire [11:0] _GEN_530 = count == 10'h18b ? _L1_wr_addr_10_T_1 : _GEN_510; // @[FSM.scala 423:28 FSM.scala 426:25]
  wire  _GEN_531 = count == 10'h18b | _GEN_511; // @[FSM.scala 423:28 FSM.scala 425:23]
  wire [11:0] _GEN_532 = count == 10'h18b ? _L1_wr_addr_11_T_1 : _GEN_512; // @[FSM.scala 423:28 FSM.scala 426:25]
  wire  _GEN_533 = count == 10'h18c | _GEN_515; // @[FSM.scala 429:28 FSM.scala 431:23]
  wire [11:0] _GEN_534 = count == 10'h18c ? _L1_wr_addr_3_T_1 : _GEN_516; // @[FSM.scala 429:28 FSM.scala 432:25]
  wire  _GEN_535 = count == 10'h18c | _GEN_517; // @[FSM.scala 429:28 FSM.scala 431:23]
  wire [11:0] _GEN_536 = count == 10'h18c ? _L1_wr_addr_4_T_1 : _GEN_518; // @[FSM.scala 429:28 FSM.scala 432:25]
  wire  _GEN_537 = count == 10'h18c | _GEN_519; // @[FSM.scala 429:28 FSM.scala 431:23]
  wire [11:0] _GEN_538 = count == 10'h18c ? _L1_wr_addr_5_T_1 : _GEN_520; // @[FSM.scala 429:28 FSM.scala 432:25]
  wire  _GEN_539 = count == 10'h18c | _GEN_521; // @[FSM.scala 429:28 FSM.scala 431:23]
  wire [11:0] _GEN_540 = count == 10'h18c ? _L1_wr_addr_6_T_1 : _GEN_522; // @[FSM.scala 429:28 FSM.scala 432:25]
  wire  _GEN_541 = count == 10'h18c | _GEN_523; // @[FSM.scala 429:28 FSM.scala 431:23]
  wire [11:0] _GEN_542 = count == 10'h18c ? _L1_wr_addr_7_T_1 : _GEN_524; // @[FSM.scala 429:28 FSM.scala 432:25]
  wire  _GEN_543 = count == 10'h18c | _GEN_525; // @[FSM.scala 429:28 FSM.scala 431:23]
  wire [11:0] _GEN_544 = count == 10'h18c ? _L1_wr_addr_8_T_1 : _GEN_526; // @[FSM.scala 429:28 FSM.scala 432:25]
  wire  _GEN_545 = count == 10'h18c | _GEN_527; // @[FSM.scala 429:28 FSM.scala 431:23]
  wire [11:0] _GEN_546 = count == 10'h18c ? _L1_wr_addr_9_T_1 : _GEN_528; // @[FSM.scala 429:28 FSM.scala 432:25]
  wire  _GEN_547 = count == 10'h18c | _GEN_529; // @[FSM.scala 429:28 FSM.scala 431:23]
  wire [11:0] _GEN_548 = count == 10'h18c ? _L1_wr_addr_10_T_1 : _GEN_530; // @[FSM.scala 429:28 FSM.scala 432:25]
  wire  _GEN_549 = count == 10'h18c | _GEN_531; // @[FSM.scala 429:28 FSM.scala 431:23]
  wire [11:0] _GEN_550 = count == 10'h18c ? _L1_wr_addr_11_T_1 : _GEN_532; // @[FSM.scala 429:28 FSM.scala 432:25]
  wire  _GEN_551 = count == 10'h18d | _GEN_535; // @[FSM.scala 435:28 FSM.scala 437:23]
  wire [11:0] _GEN_552 = count == 10'h18d ? _L1_wr_addr_4_T_1 : _GEN_536; // @[FSM.scala 435:28 FSM.scala 438:25]
  wire  _GEN_553 = count == 10'h18d | _GEN_537; // @[FSM.scala 435:28 FSM.scala 437:23]
  wire [11:0] _GEN_554 = count == 10'h18d ? _L1_wr_addr_5_T_1 : _GEN_538; // @[FSM.scala 435:28 FSM.scala 438:25]
  wire  _GEN_555 = count == 10'h18d | _GEN_539; // @[FSM.scala 435:28 FSM.scala 437:23]
  wire [11:0] _GEN_556 = count == 10'h18d ? _L1_wr_addr_6_T_1 : _GEN_540; // @[FSM.scala 435:28 FSM.scala 438:25]
  wire  _GEN_557 = count == 10'h18d | _GEN_541; // @[FSM.scala 435:28 FSM.scala 437:23]
  wire [11:0] _GEN_558 = count == 10'h18d ? _L1_wr_addr_7_T_1 : _GEN_542; // @[FSM.scala 435:28 FSM.scala 438:25]
  wire  _GEN_559 = count == 10'h18d | _GEN_543; // @[FSM.scala 435:28 FSM.scala 437:23]
  wire [11:0] _GEN_560 = count == 10'h18d ? _L1_wr_addr_8_T_1 : _GEN_544; // @[FSM.scala 435:28 FSM.scala 438:25]
  wire  _GEN_561 = count == 10'h18d | _GEN_545; // @[FSM.scala 435:28 FSM.scala 437:23]
  wire [11:0] _GEN_562 = count == 10'h18d ? _L1_wr_addr_9_T_1 : _GEN_546; // @[FSM.scala 435:28 FSM.scala 438:25]
  wire  _GEN_563 = count == 10'h18d | _GEN_547; // @[FSM.scala 435:28 FSM.scala 437:23]
  wire [11:0] _GEN_564 = count == 10'h18d ? _L1_wr_addr_10_T_1 : _GEN_548; // @[FSM.scala 435:28 FSM.scala 438:25]
  wire  _GEN_565 = count == 10'h18d | _GEN_549; // @[FSM.scala 435:28 FSM.scala 437:23]
  wire [11:0] _GEN_566 = count == 10'h18d ? _L1_wr_addr_11_T_1 : _GEN_550; // @[FSM.scala 435:28 FSM.scala 438:25]
  wire  _T_69 = count == 10'h18e; // @[FSM.scala 441:18]
  wire  _GEN_567 = count == 10'h18e | _GEN_553; // @[FSM.scala 441:28 FSM.scala 443:23]
  wire [11:0] _GEN_568 = count == 10'h18e ? _L1_wr_addr_5_T_1 : _GEN_554; // @[FSM.scala 441:28 FSM.scala 444:25]
  wire  _GEN_569 = count == 10'h18e | _GEN_555; // @[FSM.scala 441:28 FSM.scala 443:23]
  wire [11:0] _GEN_570 = count == 10'h18e ? _L1_wr_addr_6_T_1 : _GEN_556; // @[FSM.scala 441:28 FSM.scala 444:25]
  wire  _GEN_571 = count == 10'h18e | _GEN_557; // @[FSM.scala 441:28 FSM.scala 443:23]
  wire [11:0] _GEN_572 = count == 10'h18e ? _L1_wr_addr_7_T_1 : _GEN_558; // @[FSM.scala 441:28 FSM.scala 444:25]
  wire  _GEN_573 = count == 10'h18e | _GEN_559; // @[FSM.scala 441:28 FSM.scala 443:23]
  wire [11:0] _GEN_574 = count == 10'h18e ? _L1_wr_addr_8_T_1 : _GEN_560; // @[FSM.scala 441:28 FSM.scala 444:25]
  wire  _GEN_575 = count == 10'h18e | _GEN_561; // @[FSM.scala 441:28 FSM.scala 443:23]
  wire [11:0] _GEN_576 = count == 10'h18e ? _L1_wr_addr_9_T_1 : _GEN_562; // @[FSM.scala 441:28 FSM.scala 444:25]
  wire  _GEN_577 = count == 10'h18e | _GEN_563; // @[FSM.scala 441:28 FSM.scala 443:23]
  wire [11:0] _GEN_578 = count == 10'h18e ? _L1_wr_addr_10_T_1 : _GEN_564; // @[FSM.scala 441:28 FSM.scala 444:25]
  wire  _GEN_579 = count == 10'h18e | _GEN_565; // @[FSM.scala 441:28 FSM.scala 443:23]
  wire [11:0] _GEN_580 = count == 10'h18e ? _L1_wr_addr_11_T_1 : _GEN_566; // @[FSM.scala 441:28 FSM.scala 444:25]
  wire  _GEN_581 = count == 10'h18f | _GEN_569; // @[FSM.scala 447:28 FSM.scala 449:23]
  wire [11:0] _GEN_582 = count == 10'h18f ? _L1_wr_addr_6_T_1 : _GEN_570; // @[FSM.scala 447:28 FSM.scala 450:25]
  wire  _GEN_583 = count == 10'h18f | _GEN_571; // @[FSM.scala 447:28 FSM.scala 449:23]
  wire [11:0] _GEN_584 = count == 10'h18f ? _L1_wr_addr_7_T_1 : _GEN_572; // @[FSM.scala 447:28 FSM.scala 450:25]
  wire  _GEN_585 = count == 10'h18f | _GEN_573; // @[FSM.scala 447:28 FSM.scala 449:23]
  wire [11:0] _GEN_586 = count == 10'h18f ? _L1_wr_addr_8_T_1 : _GEN_574; // @[FSM.scala 447:28 FSM.scala 450:25]
  wire  _GEN_587 = count == 10'h18f | _GEN_575; // @[FSM.scala 447:28 FSM.scala 449:23]
  wire [11:0] _GEN_588 = count == 10'h18f ? _L1_wr_addr_9_T_1 : _GEN_576; // @[FSM.scala 447:28 FSM.scala 450:25]
  wire  _GEN_589 = count == 10'h18f | _GEN_577; // @[FSM.scala 447:28 FSM.scala 449:23]
  wire [11:0] _GEN_590 = count == 10'h18f ? _L1_wr_addr_10_T_1 : _GEN_578; // @[FSM.scala 447:28 FSM.scala 450:25]
  wire  _GEN_591 = count == 10'h18f | _GEN_579; // @[FSM.scala 447:28 FSM.scala 449:23]
  wire [11:0] _GEN_592 = count == 10'h18f ? _L1_wr_addr_11_T_1 : _GEN_580; // @[FSM.scala 447:28 FSM.scala 450:25]
  wire  _GEN_593 = count == 10'h190 | _GEN_583; // @[FSM.scala 453:28 FSM.scala 455:23]
  wire [11:0] _GEN_594 = count == 10'h190 ? _L1_wr_addr_7_T_1 : _GEN_584; // @[FSM.scala 453:28 FSM.scala 456:25]
  wire  _GEN_595 = count == 10'h190 | _GEN_585; // @[FSM.scala 453:28 FSM.scala 455:23]
  wire [11:0] _GEN_596 = count == 10'h190 ? _L1_wr_addr_8_T_1 : _GEN_586; // @[FSM.scala 453:28 FSM.scala 456:25]
  wire  _GEN_597 = count == 10'h190 | _GEN_587; // @[FSM.scala 453:28 FSM.scala 455:23]
  wire [11:0] _GEN_598 = count == 10'h190 ? _L1_wr_addr_9_T_1 : _GEN_588; // @[FSM.scala 453:28 FSM.scala 456:25]
  wire  _GEN_599 = count == 10'h190 | _GEN_589; // @[FSM.scala 453:28 FSM.scala 455:23]
  wire [11:0] _GEN_600 = count == 10'h190 ? _L1_wr_addr_10_T_1 : _GEN_590; // @[FSM.scala 453:28 FSM.scala 456:25]
  wire  _GEN_601 = count == 10'h190 | _GEN_591; // @[FSM.scala 453:28 FSM.scala 455:23]
  wire [11:0] _GEN_602 = count == 10'h190 ? _L1_wr_addr_11_T_1 : _GEN_592; // @[FSM.scala 453:28 FSM.scala 456:25]
  wire  _GEN_603 = count == 10'h191 | _GEN_595; // @[FSM.scala 459:28 FSM.scala 461:23]
  wire [11:0] _GEN_604 = count == 10'h191 ? _L1_wr_addr_8_T_1 : _GEN_596; // @[FSM.scala 459:28 FSM.scala 462:25]
  wire  _GEN_605 = count == 10'h191 | _GEN_597; // @[FSM.scala 459:28 FSM.scala 461:23]
  wire [11:0] _GEN_606 = count == 10'h191 ? _L1_wr_addr_9_T_1 : _GEN_598; // @[FSM.scala 459:28 FSM.scala 462:25]
  wire  _GEN_607 = count == 10'h191 | _GEN_599; // @[FSM.scala 459:28 FSM.scala 461:23]
  wire [11:0] _GEN_608 = count == 10'h191 ? _L1_wr_addr_10_T_1 : _GEN_600; // @[FSM.scala 459:28 FSM.scala 462:25]
  wire  _GEN_609 = count == 10'h191 | _GEN_601; // @[FSM.scala 459:28 FSM.scala 461:23]
  wire [11:0] _GEN_610 = count == 10'h191 ? _L1_wr_addr_11_T_1 : _GEN_602; // @[FSM.scala 459:28 FSM.scala 462:25]
  wire  _GEN_611 = count == 10'h192 | _GEN_605; // @[FSM.scala 465:28 FSM.scala 467:23]
  wire [11:0] _GEN_612 = count == 10'h192 ? _L1_wr_addr_9_T_1 : _GEN_606; // @[FSM.scala 465:28 FSM.scala 468:25]
  wire  _GEN_613 = count == 10'h192 | _GEN_607; // @[FSM.scala 465:28 FSM.scala 467:23]
  wire [11:0] _GEN_614 = count == 10'h192 ? _L1_wr_addr_10_T_1 : _GEN_608; // @[FSM.scala 465:28 FSM.scala 468:25]
  wire  _GEN_615 = count == 10'h192 | _GEN_609; // @[FSM.scala 465:28 FSM.scala 467:23]
  wire [11:0] _GEN_616 = count == 10'h192 ? _L1_wr_addr_11_T_1 : _GEN_610; // @[FSM.scala 465:28 FSM.scala 468:25]
  wire  _GEN_617 = count == 10'h193 | _GEN_613; // @[FSM.scala 471:28 FSM.scala 473:23]
  wire [11:0] _GEN_618 = count == 10'h193 ? _L1_wr_addr_10_T_1 : _GEN_614; // @[FSM.scala 471:28 FSM.scala 474:25]
  wire  _GEN_619 = count == 10'h193 | _GEN_615; // @[FSM.scala 471:28 FSM.scala 473:23]
  wire [11:0] _GEN_620 = count == 10'h193 ? _L1_wr_addr_11_T_1 : _GEN_616; // @[FSM.scala 471:28 FSM.scala 474:25]
  wire  _GEN_621 = count == 10'h194 | _GEN_619; // @[FSM.scala 477:28 FSM.scala 479:23]
  wire [11:0] _GEN_622 = count == 10'h194 ? _L1_wr_addr_11_T_1 : _GEN_620; // @[FSM.scala 477:28 FSM.scala 480:25]
  wire  _GEN_623 = count == 10'h195 ? 1'h0 : _GEN_467; // @[FSM.scala 484:28 FSM.scala 486:23]
  wire  _GEN_624 = count == 10'h195 ? 1'h0 : _GEN_491; // @[FSM.scala 484:28 FSM.scala 486:23]
  wire  _GEN_625 = count == 10'h195 ? 1'h0 : _GEN_513; // @[FSM.scala 484:28 FSM.scala 486:23]
  wire  _GEN_626 = count == 10'h195 ? 1'h0 : _GEN_533; // @[FSM.scala 484:28 FSM.scala 486:23]
  wire  _GEN_627 = count == 10'h195 ? 1'h0 : _GEN_551; // @[FSM.scala 484:28 FSM.scala 486:23]
  wire  _GEN_628 = count == 10'h195 ? 1'h0 : _GEN_567; // @[FSM.scala 484:28 FSM.scala 486:23]
  wire  _GEN_629 = count == 10'h195 ? 1'h0 : _GEN_581; // @[FSM.scala 484:28 FSM.scala 486:23]
  wire  _GEN_630 = count == 10'h195 ? 1'h0 : _GEN_593; // @[FSM.scala 484:28 FSM.scala 486:23]
  wire  _GEN_631 = count == 10'h195 ? 1'h0 : _GEN_603; // @[FSM.scala 484:28 FSM.scala 486:23]
  wire  _GEN_632 = count == 10'h195 ? 1'h0 : _GEN_611; // @[FSM.scala 484:28 FSM.scala 486:23]
  wire  _GEN_633 = count == 10'h195 ? 1'h0 : _GEN_617; // @[FSM.scala 484:28 FSM.scala 486:23]
  wire  _GEN_634 = count == 10'h195 ? 1'h0 : _GEN_621; // @[FSM.scala 484:28 FSM.scala 486:23]
  wire [9:0] _GEN_635 = count == 10'h195 ? 10'h0 : _GEN_234; // @[FSM.scala 484:28 FSM.scala 488:15]
  wire [6:0] _GEN_636 = count == 10'h195 ? 7'h0 : _count1_T_1; // @[FSM.scala 484:28 FSM.scala 489:16]
  wire [2:0] _GEN_638 = count == 10'h195 ? 3'h4 : state; // @[FSM.scala 484:28 FSM.scala 491:15 FSM.scala 159:22]
  wire  _T_77 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire [9:0] _GEN_639 = count != 10'h12 ? _count_T_1 : count; // @[FSM.scala 498:29 FSM.scala 499:17 FSM.scala 161:22]
  wire [2:0] _GEN_640 = _T_3 ? 3'h3 : PEArray_ctrl_2_control; // @[FSM.scala 502:28 FSM.scala 504:35 FSM.scala 64:28]
  wire [9:0] _GEN_642 = _T_3 ? 10'hf : PEArray_ctrl_2_count; // @[FSM.scala 502:28 FSM.scala 506:33 FSM.scala 64:28]
  wire [5:0] _GEN_643 = _T_3 ? 6'hf : PEArray_ctrl_2_L0index; // @[FSM.scala 502:28 FSM.scala 507:35 FSM.scala 64:28]
  wire [1:0] _GEN_644 = _T_3 ? 2'h1 : PE_above_data_ctrl; // @[FSM.scala 502:28 FSM.scala 509:30 FSM.scala 74:35]
  wire [11:0] _GEN_646 = _T_5 ? 12'h0 : PEArray_ctrl_0_mask; // @[FSM.scala 512:28 FSM.scala 514:34 FSM.scala 64:28]
  wire [11:0] _GEN_647 = _T_5 ? 12'h0 : PEArray_ctrl_1_mask; // @[FSM.scala 512:28 FSM.scala 514:34 FSM.scala 64:28]
  wire [2:0] _GEN_649 = _T_48 ? 3'h0 : Ht_to_PE_control; // @[FSM.scala 517:28 FSM.scala 518:28 FSM.scala 77:36]
  wire  _T_85 = count >= 10'h3 & count <= 10'h7; // @[FSM.scala 521:29]
  wire [2:0] _Ht_to_PE_control_T_1 = Ht_to_PE_control + 3'h1; // @[FSM.scala 522:48]
  wire [2:0] _GEN_650 = count >= 10'h3 & count <= 10'h7 ? _Ht_to_PE_control_T_1 : _GEN_649; // @[FSM.scala 521:47 FSM.scala 522:28]
  wire [1:0] _GEN_651 = _T_53 ? 2'h0 : _GEN_644; // @[FSM.scala 525:28 FSM.scala 526:30]
  wire [11:0] _GEN_652 = _T_53 ? 12'h0 : L1_rd_addr_0; // @[FSM.scala 525:28 FSM.scala 528:27 FSM.scala 60:28]
  wire [11:0] _GEN_653 = _T_53 ? 12'h0 : L1_rd_addr_1; // @[FSM.scala 525:28 FSM.scala 528:27 FSM.scala 60:28]
  wire [11:0] _GEN_654 = _T_53 ? 12'h0 : L1_rd_addr_2; // @[FSM.scala 525:28 FSM.scala 528:27 FSM.scala 60:28]
  wire [11:0] _GEN_655 = _T_53 ? 12'h0 : L1_rd_addr_3; // @[FSM.scala 525:28 FSM.scala 528:27 FSM.scala 60:28]
  wire [11:0] _GEN_656 = _T_53 ? 12'h0 : L1_rd_addr_4; // @[FSM.scala 525:28 FSM.scala 528:27 FSM.scala 60:28]
  wire [11:0] _GEN_657 = _T_53 ? 12'h0 : L1_rd_addr_5; // @[FSM.scala 525:28 FSM.scala 528:27 FSM.scala 60:28]
  wire [11:0] _GEN_658 = _T_53 ? 12'h0 : L1_rd_addr_6; // @[FSM.scala 525:28 FSM.scala 528:27 FSM.scala 60:28]
  wire [11:0] _GEN_659 = _T_53 ? 12'h0 : L1_rd_addr_7; // @[FSM.scala 525:28 FSM.scala 528:27 FSM.scala 60:28]
  wire [11:0] _GEN_660 = _T_53 ? 12'h0 : L1_rd_addr_8; // @[FSM.scala 525:28 FSM.scala 528:27 FSM.scala 60:28]
  wire [11:0] _GEN_661 = _T_53 ? 12'h0 : L1_rd_addr_9; // @[FSM.scala 525:28 FSM.scala 528:27 FSM.scala 60:28]
  wire [11:0] _GEN_662 = _T_53 ? 12'h0 : L1_rd_addr_10; // @[FSM.scala 525:28 FSM.scala 528:27 FSM.scala 60:28]
  wire [11:0] _GEN_663 = _T_53 ? 12'h0 : L1_rd_addr_11; // @[FSM.scala 525:28 FSM.scala 528:27 FSM.scala 60:28]
  wire [11:0] _GEN_664 = count >= 10'h8 & count <= 10'he ? _L1_rd_addr_0_T_1 : _GEN_652; // @[FSM.scala 532:48 FSM.scala 534:27]
  wire [11:0] _GEN_665 = count >= 10'h8 & count <= 10'he ? _L1_rd_addr_1_T_1 : _GEN_653; // @[FSM.scala 532:48 FSM.scala 534:27]
  wire [11:0] _GEN_666 = count >= 10'h8 & count <= 10'he ? _L1_rd_addr_2_T_1 : _GEN_654; // @[FSM.scala 532:48 FSM.scala 534:27]
  wire [11:0] _GEN_667 = count >= 10'h8 & count <= 10'he ? _L1_rd_addr_3_T_1 : _GEN_655; // @[FSM.scala 532:48 FSM.scala 534:27]
  wire [11:0] _GEN_668 = count >= 10'h8 & count <= 10'he ? _L1_rd_addr_4_T_1 : _GEN_656; // @[FSM.scala 532:48 FSM.scala 534:27]
  wire [11:0] _GEN_669 = count >= 10'h8 & count <= 10'he ? _L1_rd_addr_5_T_1 : _GEN_657; // @[FSM.scala 532:48 FSM.scala 534:27]
  wire [11:0] _GEN_670 = count >= 10'h8 & count <= 10'he ? _L1_rd_addr_6_T_1 : _GEN_658; // @[FSM.scala 532:48 FSM.scala 534:27]
  wire [11:0] _GEN_671 = count >= 10'h8 & count <= 10'he ? _L1_rd_addr_7_T_1 : _GEN_659; // @[FSM.scala 532:48 FSM.scala 534:27]
  wire [11:0] _GEN_672 = count >= 10'h8 & count <= 10'he ? _L1_rd_addr_8_T_1 : _GEN_660; // @[FSM.scala 532:48 FSM.scala 534:27]
  wire [11:0] _GEN_673 = count >= 10'h8 & count <= 10'he ? _L1_rd_addr_9_T_1 : _GEN_661; // @[FSM.scala 532:48 FSM.scala 534:27]
  wire [11:0] _GEN_674 = count >= 10'h8 & count <= 10'he ? _L1_rd_addr_10_T_1 : _GEN_662; // @[FSM.scala 532:48 FSM.scala 534:27]
  wire [11:0] _GEN_675 = count >= 10'h8 & count <= 10'he ? _L1_rd_addr_11_T_1 : _GEN_663; // @[FSM.scala 532:48 FSM.scala 534:27]
  wire [9:0] _GEN_676 = count == 10'h12 ? 10'h0 : _GEN_639; // @[FSM.scala 537:29 FSM.scala 538:17]
  wire [3:0] _GEN_677 = count == 10'h12 ? 4'h1 : gru_state; // @[FSM.scala 537:29 FSM.scala 539:21 FSM.scala 160:26]
  wire [9:0] _GEN_678 = gru_state == 4'h0 ? _GEN_676 : count; // @[FSM.scala 497:30 FSM.scala 161:22]
  wire [2:0] _GEN_679 = gru_state == 4'h0 ? _GEN_640 : PEArray_ctrl_2_control; // @[FSM.scala 497:30 FSM.scala 64:28]
  wire [11:0] _GEN_680 = gru_state == 4'h0 ? _GEN_108 : PEArray_ctrl_2_mask; // @[FSM.scala 497:30 FSM.scala 64:28]
  wire [9:0] _GEN_681 = gru_state == 4'h0 ? _GEN_642 : PEArray_ctrl_2_count; // @[FSM.scala 497:30 FSM.scala 64:28]
  wire [5:0] _GEN_682 = gru_state == 4'h0 ? _GEN_643 : PEArray_ctrl_2_L0index; // @[FSM.scala 497:30 FSM.scala 64:28]
  wire [1:0] _GEN_683 = gru_state == 4'h0 ? _GEN_651 : PE_above_data_ctrl; // @[FSM.scala 497:30 FSM.scala 74:35]
  wire [3:0] _GEN_684 = gru_state == 4'h0 ? _GEN_105 : PE_rd_data_mux; // @[FSM.scala 497:30 FSM.scala 61:32]
  wire [11:0] _GEN_685 = gru_state == 4'h0 ? _GEN_646 : PEArray_ctrl_0_mask; // @[FSM.scala 497:30 FSM.scala 64:28]
  wire [11:0] _GEN_686 = gru_state == 4'h0 ? _GEN_647 : PEArray_ctrl_1_mask; // @[FSM.scala 497:30 FSM.scala 64:28]
  wire [2:0] _GEN_687 = gru_state == 4'h0 ? _GEN_650 : Ht_to_PE_control; // @[FSM.scala 497:30 FSM.scala 77:36]
  wire [11:0] _GEN_688 = gru_state == 4'h0 ? _GEN_664 : L1_rd_addr_0; // @[FSM.scala 497:30 FSM.scala 60:28]
  wire [11:0] _GEN_689 = gru_state == 4'h0 ? _GEN_665 : L1_rd_addr_1; // @[FSM.scala 497:30 FSM.scala 60:28]
  wire [11:0] _GEN_690 = gru_state == 4'h0 ? _GEN_666 : L1_rd_addr_2; // @[FSM.scala 497:30 FSM.scala 60:28]
  wire [11:0] _GEN_691 = gru_state == 4'h0 ? _GEN_667 : L1_rd_addr_3; // @[FSM.scala 497:30 FSM.scala 60:28]
  wire [11:0] _GEN_692 = gru_state == 4'h0 ? _GEN_668 : L1_rd_addr_4; // @[FSM.scala 497:30 FSM.scala 60:28]
  wire [11:0] _GEN_693 = gru_state == 4'h0 ? _GEN_669 : L1_rd_addr_5; // @[FSM.scala 497:30 FSM.scala 60:28]
  wire [11:0] _GEN_694 = gru_state == 4'h0 ? _GEN_670 : L1_rd_addr_6; // @[FSM.scala 497:30 FSM.scala 60:28]
  wire [11:0] _GEN_695 = gru_state == 4'h0 ? _GEN_671 : L1_rd_addr_7; // @[FSM.scala 497:30 FSM.scala 60:28]
  wire [11:0] _GEN_696 = gru_state == 4'h0 ? _GEN_672 : L1_rd_addr_8; // @[FSM.scala 497:30 FSM.scala 60:28]
  wire [11:0] _GEN_697 = gru_state == 4'h0 ? _GEN_673 : L1_rd_addr_9; // @[FSM.scala 497:30 FSM.scala 60:28]
  wire [11:0] _GEN_698 = gru_state == 4'h0 ? _GEN_674 : L1_rd_addr_10; // @[FSM.scala 497:30 FSM.scala 60:28]
  wire [11:0] _GEN_699 = gru_state == 4'h0 ? _GEN_675 : L1_rd_addr_11; // @[FSM.scala 497:30 FSM.scala 60:28]
  wire [3:0] _GEN_700 = gru_state == 4'h0 ? _GEN_677 : gru_state; // @[FSM.scala 497:30 FSM.scala 160:26]
  wire  _T_92 = count != 10'h38e; // @[FSM.scala 544:20]
  wire [9:0] _GEN_701 = count != 10'h38e ? _count_T_1 : _GEN_678; // @[FSM.scala 544:30 FSM.scala 545:17]
  wire [6:0] _GEN_702 = count1 != 7'h3f ? _count1_T_1 : 7'h0; // @[FSM.scala 548:30 FSM.scala 549:18 FSM.scala 551:18]
  wire [2:0] _GEN_703 = _T_3 ? 3'h4 : _GEN_679; // @[FSM.scala 554:28 FSM.scala 556:35]
  wire [9:0] _GEN_704 = _T_3 ? 10'h37f : _GEN_681; // @[FSM.scala 554:28 FSM.scala 557:33]
  wire [5:0] _GEN_705 = _T_3 ? 6'hf : _GEN_682; // @[FSM.scala 554:28 FSM.scala 558:35]
  wire [11:0] _GEN_706 = _T_3 ? 12'h800 : _GEN_680; // @[FSM.scala 554:28 FSM.scala 559:32]
  wire [7:0] _GEN_707 = _T_3 ? 8'h40 : PEArray_ctrl_2_gru_out_width; // @[FSM.scala 554:28 FSM.scala 560:41 FSM.scala 64:28]
  wire [11:0] _GEN_708 = _T_3 ? 12'h1f4 : _GEN_688; // @[FSM.scala 554:28 FSM.scala 564:27]
  wire [11:0] _GEN_709 = _T_3 ? 12'h1f4 : _GEN_689; // @[FSM.scala 554:28 FSM.scala 564:27]
  wire [11:0] _GEN_710 = _T_3 ? 12'h1f4 : _GEN_690; // @[FSM.scala 554:28 FSM.scala 564:27]
  wire [11:0] _GEN_711 = _T_3 ? 12'h1f4 : _GEN_691; // @[FSM.scala 554:28 FSM.scala 564:27]
  wire [11:0] _GEN_712 = _T_3 ? 12'h1f4 : _GEN_692; // @[FSM.scala 554:28 FSM.scala 564:27]
  wire [11:0] _GEN_713 = _T_3 ? 12'h1f4 : _GEN_693; // @[FSM.scala 554:28 FSM.scala 564:27]
  wire [11:0] _GEN_714 = _T_3 ? 12'h1f4 : _GEN_694; // @[FSM.scala 554:28 FSM.scala 564:27]
  wire [11:0] _GEN_715 = _T_3 ? 12'h1f4 : _GEN_695; // @[FSM.scala 554:28 FSM.scala 564:27]
  wire [11:0] _GEN_716 = _T_3 ? 12'h1f4 : _GEN_696; // @[FSM.scala 554:28 FSM.scala 564:27]
  wire [11:0] _GEN_717 = _T_3 ? 12'h1f4 : _GEN_697; // @[FSM.scala 554:28 FSM.scala 564:27]
  wire [11:0] _GEN_718 = _T_3 ? 12'h1f4 : _GEN_698; // @[FSM.scala 554:28 FSM.scala 564:27]
  wire [11:0] _GEN_719 = _T_3 ? 12'h1f4 : _GEN_699; // @[FSM.scala 554:28 FSM.scala 564:27]
  wire [1:0] _GEN_720 = _T_3 ? 2'h0 : _GEN_683; // @[FSM.scala 554:28 FSM.scala 566:30]
  wire [3:0] _GEN_721 = _T_3 ? 4'h0 : _GEN_684; // @[FSM.scala 554:28 FSM.scala 567:26]
  wire [5:0] _GEN_722 = _T_3 ? 6'h0 : Zt_wrAddr; // @[FSM.scala 554:28 FSM.scala 570:21 FSM.scala 83:36]
  wire [1:0] _GEN_723 = _T_3 ? 2'h1 : BN_Unit_ctrl; // @[FSM.scala 554:28 FSM.scala 571:24 FSM.scala 69:28]
  wire [1:0] _GEN_724 = _T_3 ? 2'h1 : Activation_ctrl; // @[FSM.scala 554:28 FSM.scala 572:27 FSM.scala 75:32]
  wire [2:0] _GEN_725 = _T_39 ? 3'h4 : _GEN_703; // @[FSM.scala 576:48 FSM.scala 577:35]
  wire [9:0] _GEN_726 = _T_39 ? 10'h37f : _GEN_704; // @[FSM.scala 576:48 FSM.scala 578:33]
  wire [5:0] _GEN_727 = _T_39 ? 6'hf : _GEN_705; // @[FSM.scala 576:48 FSM.scala 579:35]
  wire [11:0] _GEN_728 = _T_39 ? {{1'd0}, PEArray_ctrl_2_mask[11:1]} : _GEN_706; // @[FSM.scala 576:48 FSM.scala 580:32]
  wire [7:0] _GEN_729 = _T_39 ? 8'h40 : _GEN_707; // @[FSM.scala 576:48 FSM.scala 581:41]
  wire [11:0] _GEN_730 = _T_40 ? 12'h0 : _GEN_685; // @[FSM.scala 583:29 FSM.scala 585:34]
  wire [11:0] _GEN_731 = _T_40 ? 12'h0 : _GEN_686; // @[FSM.scala 583:29 FSM.scala 585:34]
  wire [11:0] _GEN_732 = _T_40 ? 12'h0 : _GEN_728; // @[FSM.scala 583:29 FSM.scala 585:34]
  wire [11:0] _GEN_733 = _T_5 ? _L1_rd_addr_0_T_1 : _GEN_708; // @[FSM.scala 590:28 FSM.scala 592:27]
  wire [11:0] _GEN_734 = _T_48 ? _L1_rd_addr_0_T_1 : _GEN_733; // @[FSM.scala 595:28 FSM.scala 597:27]
  wire [11:0] _GEN_735 = _T_48 ? _L1_rd_addr_1_T_1 : _GEN_709; // @[FSM.scala 595:28 FSM.scala 597:27]
  wire [11:0] _GEN_736 = _T_49 ? _L1_rd_addr_0_T_1 : _GEN_734; // @[FSM.scala 600:28 FSM.scala 602:27]
  wire [11:0] _GEN_737 = _T_49 ? _L1_rd_addr_1_T_1 : _GEN_735; // @[FSM.scala 600:28 FSM.scala 602:27]
  wire [11:0] _GEN_738 = _T_49 ? _L1_rd_addr_2_T_1 : _GEN_710; // @[FSM.scala 600:28 FSM.scala 602:27]
  wire [11:0] _GEN_739 = _T_21 ? _L1_rd_addr_0_T_1 : _GEN_736; // @[FSM.scala 605:28 FSM.scala 607:27]
  wire [11:0] _GEN_740 = _T_21 ? _L1_rd_addr_1_T_1 : _GEN_737; // @[FSM.scala 605:28 FSM.scala 607:27]
  wire [11:0] _GEN_741 = _T_21 ? _L1_rd_addr_2_T_1 : _GEN_738; // @[FSM.scala 605:28 FSM.scala 607:27]
  wire [11:0] _GEN_742 = _T_21 ? _L1_rd_addr_3_T_1 : _GEN_711; // @[FSM.scala 605:28 FSM.scala 607:27]
  wire [11:0] _GEN_743 = _T_51 ? _L1_rd_addr_0_T_1 : _GEN_739; // @[FSM.scala 610:28 FSM.scala 612:27]
  wire [11:0] _GEN_744 = _T_51 ? _L1_rd_addr_1_T_1 : _GEN_740; // @[FSM.scala 610:28 FSM.scala 612:27]
  wire [11:0] _GEN_745 = _T_51 ? _L1_rd_addr_2_T_1 : _GEN_741; // @[FSM.scala 610:28 FSM.scala 612:27]
  wire [11:0] _GEN_746 = _T_51 ? _L1_rd_addr_3_T_1 : _GEN_742; // @[FSM.scala 610:28 FSM.scala 612:27]
  wire [11:0] _GEN_747 = _T_51 ? _L1_rd_addr_4_T_1 : _GEN_712; // @[FSM.scala 610:28 FSM.scala 612:27]
  wire [11:0] _GEN_748 = _T_52 ? _L1_rd_addr_0_T_1 : _GEN_743; // @[FSM.scala 615:28 FSM.scala 617:27]
  wire [11:0] _GEN_749 = _T_52 ? _L1_rd_addr_1_T_1 : _GEN_744; // @[FSM.scala 615:28 FSM.scala 617:27]
  wire [11:0] _GEN_750 = _T_52 ? _L1_rd_addr_2_T_1 : _GEN_745; // @[FSM.scala 615:28 FSM.scala 617:27]
  wire [11:0] _GEN_751 = _T_52 ? _L1_rd_addr_3_T_1 : _GEN_746; // @[FSM.scala 615:28 FSM.scala 617:27]
  wire [11:0] _GEN_752 = _T_52 ? _L1_rd_addr_4_T_1 : _GEN_747; // @[FSM.scala 615:28 FSM.scala 617:27]
  wire [11:0] _GEN_753 = _T_52 ? _L1_rd_addr_5_T_1 : _GEN_713; // @[FSM.scala 615:28 FSM.scala 617:27]
  wire [11:0] _GEN_754 = _T_53 ? _L1_rd_addr_0_T_1 : _GEN_748; // @[FSM.scala 620:28 FSM.scala 622:27]
  wire [11:0] _GEN_755 = _T_53 ? _L1_rd_addr_1_T_1 : _GEN_749; // @[FSM.scala 620:28 FSM.scala 622:27]
  wire [11:0] _GEN_756 = _T_53 ? _L1_rd_addr_2_T_1 : _GEN_750; // @[FSM.scala 620:28 FSM.scala 622:27]
  wire [11:0] _GEN_757 = _T_53 ? _L1_rd_addr_3_T_1 : _GEN_751; // @[FSM.scala 620:28 FSM.scala 622:27]
  wire [11:0] _GEN_758 = _T_53 ? _L1_rd_addr_4_T_1 : _GEN_752; // @[FSM.scala 620:28 FSM.scala 622:27]
  wire [11:0] _GEN_759 = _T_53 ? _L1_rd_addr_5_T_1 : _GEN_753; // @[FSM.scala 620:28 FSM.scala 622:27]
  wire [11:0] _GEN_760 = _T_53 ? _L1_rd_addr_6_T_1 : _GEN_714; // @[FSM.scala 620:28 FSM.scala 622:27]
  wire [11:0] _GEN_761 = _T_54 ? _L1_rd_addr_0_T_1 : _GEN_754; // @[FSM.scala 625:28 FSM.scala 627:27]
  wire [11:0] _GEN_762 = _T_54 ? _L1_rd_addr_1_T_1 : _GEN_755; // @[FSM.scala 625:28 FSM.scala 627:27]
  wire [11:0] _GEN_763 = _T_54 ? _L1_rd_addr_2_T_1 : _GEN_756; // @[FSM.scala 625:28 FSM.scala 627:27]
  wire [11:0] _GEN_764 = _T_54 ? _L1_rd_addr_3_T_1 : _GEN_757; // @[FSM.scala 625:28 FSM.scala 627:27]
  wire [11:0] _GEN_765 = _T_54 ? _L1_rd_addr_4_T_1 : _GEN_758; // @[FSM.scala 625:28 FSM.scala 627:27]
  wire [11:0] _GEN_766 = _T_54 ? _L1_rd_addr_5_T_1 : _GEN_759; // @[FSM.scala 625:28 FSM.scala 627:27]
  wire [11:0] _GEN_767 = _T_54 ? _L1_rd_addr_6_T_1 : _GEN_760; // @[FSM.scala 625:28 FSM.scala 627:27]
  wire [11:0] _GEN_768 = _T_54 ? _L1_rd_addr_7_T_1 : _GEN_715; // @[FSM.scala 625:28 FSM.scala 627:27]
  wire [11:0] _GEN_769 = _T_55 ? _L1_rd_addr_0_T_1 : _GEN_761; // @[FSM.scala 630:28 FSM.scala 632:27]
  wire [11:0] _GEN_770 = _T_55 ? _L1_rd_addr_1_T_1 : _GEN_762; // @[FSM.scala 630:28 FSM.scala 632:27]
  wire [11:0] _GEN_771 = _T_55 ? _L1_rd_addr_2_T_1 : _GEN_763; // @[FSM.scala 630:28 FSM.scala 632:27]
  wire [11:0] _GEN_772 = _T_55 ? _L1_rd_addr_3_T_1 : _GEN_764; // @[FSM.scala 630:28 FSM.scala 632:27]
  wire [11:0] _GEN_773 = _T_55 ? _L1_rd_addr_4_T_1 : _GEN_765; // @[FSM.scala 630:28 FSM.scala 632:27]
  wire [11:0] _GEN_774 = _T_55 ? _L1_rd_addr_5_T_1 : _GEN_766; // @[FSM.scala 630:28 FSM.scala 632:27]
  wire [11:0] _GEN_775 = _T_55 ? _L1_rd_addr_6_T_1 : _GEN_767; // @[FSM.scala 630:28 FSM.scala 632:27]
  wire [11:0] _GEN_776 = _T_55 ? _L1_rd_addr_7_T_1 : _GEN_768; // @[FSM.scala 630:28 FSM.scala 632:27]
  wire [11:0] _GEN_777 = _T_55 ? _L1_rd_addr_8_T_1 : _GEN_716; // @[FSM.scala 630:28 FSM.scala 632:27]
  wire [11:0] _GEN_778 = _T_56 ? _L1_rd_addr_0_T_1 : _GEN_769; // @[FSM.scala 635:29 FSM.scala 637:27]
  wire [11:0] _GEN_779 = _T_56 ? _L1_rd_addr_1_T_1 : _GEN_770; // @[FSM.scala 635:29 FSM.scala 637:27]
  wire [11:0] _GEN_780 = _T_56 ? _L1_rd_addr_2_T_1 : _GEN_771; // @[FSM.scala 635:29 FSM.scala 637:27]
  wire [11:0] _GEN_781 = _T_56 ? _L1_rd_addr_3_T_1 : _GEN_772; // @[FSM.scala 635:29 FSM.scala 637:27]
  wire [11:0] _GEN_782 = _T_56 ? _L1_rd_addr_4_T_1 : _GEN_773; // @[FSM.scala 635:29 FSM.scala 637:27]
  wire [11:0] _GEN_783 = _T_56 ? _L1_rd_addr_5_T_1 : _GEN_774; // @[FSM.scala 635:29 FSM.scala 637:27]
  wire [11:0] _GEN_784 = _T_56 ? _L1_rd_addr_6_T_1 : _GEN_775; // @[FSM.scala 635:29 FSM.scala 637:27]
  wire [11:0] _GEN_785 = _T_56 ? _L1_rd_addr_7_T_1 : _GEN_776; // @[FSM.scala 635:29 FSM.scala 637:27]
  wire [11:0] _GEN_786 = _T_56 ? _L1_rd_addr_8_T_1 : _GEN_777; // @[FSM.scala 635:29 FSM.scala 637:27]
  wire [11:0] _GEN_787 = _T_56 ? _L1_rd_addr_9_T_1 : _GEN_717; // @[FSM.scala 635:29 FSM.scala 637:27]
  wire [11:0] _GEN_788 = _T_57 ? _L1_rd_addr_0_T_1 : _GEN_778; // @[FSM.scala 640:29 FSM.scala 642:27]
  wire [11:0] _GEN_789 = _T_57 ? _L1_rd_addr_1_T_1 : _GEN_779; // @[FSM.scala 640:29 FSM.scala 642:27]
  wire [11:0] _GEN_790 = _T_57 ? _L1_rd_addr_2_T_1 : _GEN_780; // @[FSM.scala 640:29 FSM.scala 642:27]
  wire [11:0] _GEN_791 = _T_57 ? _L1_rd_addr_3_T_1 : _GEN_781; // @[FSM.scala 640:29 FSM.scala 642:27]
  wire [11:0] _GEN_792 = _T_57 ? _L1_rd_addr_4_T_1 : _GEN_782; // @[FSM.scala 640:29 FSM.scala 642:27]
  wire [11:0] _GEN_793 = _T_57 ? _L1_rd_addr_5_T_1 : _GEN_783; // @[FSM.scala 640:29 FSM.scala 642:27]
  wire [11:0] _GEN_794 = _T_57 ? _L1_rd_addr_6_T_1 : _GEN_784; // @[FSM.scala 640:29 FSM.scala 642:27]
  wire [11:0] _GEN_795 = _T_57 ? _L1_rd_addr_7_T_1 : _GEN_785; // @[FSM.scala 640:29 FSM.scala 642:27]
  wire [11:0] _GEN_796 = _T_57 ? _L1_rd_addr_8_T_1 : _GEN_786; // @[FSM.scala 640:29 FSM.scala 642:27]
  wire [11:0] _GEN_797 = _T_57 ? _L1_rd_addr_9_T_1 : _GEN_787; // @[FSM.scala 640:29 FSM.scala 642:27]
  wire [11:0] _GEN_798 = _T_57 ? _L1_rd_addr_10_T_1 : _GEN_718; // @[FSM.scala 640:29 FSM.scala 642:27]
  wire  _T_110 = count >= 10'hc; // @[FSM.scala 645:21]
  wire  _T_112 = count >= 10'hc & count <= 10'h37f; // @[FSM.scala 645:30]
  wire [11:0] _GEN_799 = count >= 10'hc & count <= 10'h37f ? _L1_rd_addr_0_T_1 : _GEN_788; // @[FSM.scala 645:50 FSM.scala 647:27]
  wire [11:0] _GEN_800 = count >= 10'hc & count <= 10'h37f ? _L1_rd_addr_1_T_1 : _GEN_789; // @[FSM.scala 645:50 FSM.scala 647:27]
  wire [11:0] _GEN_801 = count >= 10'hc & count <= 10'h37f ? _L1_rd_addr_2_T_1 : _GEN_790; // @[FSM.scala 645:50 FSM.scala 647:27]
  wire [11:0] _GEN_802 = count >= 10'hc & count <= 10'h37f ? _L1_rd_addr_3_T_1 : _GEN_791; // @[FSM.scala 645:50 FSM.scala 647:27]
  wire [11:0] _GEN_803 = count >= 10'hc & count <= 10'h37f ? _L1_rd_addr_4_T_1 : _GEN_792; // @[FSM.scala 645:50 FSM.scala 647:27]
  wire [11:0] _GEN_804 = count >= 10'hc & count <= 10'h37f ? _L1_rd_addr_5_T_1 : _GEN_793; // @[FSM.scala 645:50 FSM.scala 647:27]
  wire [11:0] _GEN_805 = count >= 10'hc & count <= 10'h37f ? _L1_rd_addr_6_T_1 : _GEN_794; // @[FSM.scala 645:50 FSM.scala 647:27]
  wire [11:0] _GEN_806 = count >= 10'hc & count <= 10'h37f ? _L1_rd_addr_7_T_1 : _GEN_795; // @[FSM.scala 645:50 FSM.scala 647:27]
  wire [11:0] _GEN_807 = count >= 10'hc & count <= 10'h37f ? _L1_rd_addr_8_T_1 : _GEN_796; // @[FSM.scala 645:50 FSM.scala 647:27]
  wire [11:0] _GEN_808 = count >= 10'hc & count <= 10'h37f ? _L1_rd_addr_9_T_1 : _GEN_797; // @[FSM.scala 645:50 FSM.scala 647:27]
  wire [11:0] _GEN_809 = count >= 10'hc & count <= 10'h37f ? _L1_rd_addr_10_T_1 : _GEN_798; // @[FSM.scala 645:50 FSM.scala 647:27]
  wire [11:0] _GEN_810 = count >= 10'hc & count <= 10'h37f ? _L1_rd_addr_11_T_1 : _GEN_719; // @[FSM.scala 645:50 FSM.scala 647:27]
  wire  _T_113 = count == 10'h380; // @[FSM.scala 650:20]
  wire [11:0] _GEN_811 = count == 10'h380 ? _L1_rd_addr_1_T_1 : _GEN_800; // @[FSM.scala 650:30 FSM.scala 652:27]
  wire [11:0] _GEN_812 = count == 10'h380 ? _L1_rd_addr_2_T_1 : _GEN_801; // @[FSM.scala 650:30 FSM.scala 652:27]
  wire [11:0] _GEN_813 = count == 10'h380 ? _L1_rd_addr_3_T_1 : _GEN_802; // @[FSM.scala 650:30 FSM.scala 652:27]
  wire [11:0] _GEN_814 = count == 10'h380 ? _L1_rd_addr_4_T_1 : _GEN_803; // @[FSM.scala 650:30 FSM.scala 652:27]
  wire [11:0] _GEN_815 = count == 10'h380 ? _L1_rd_addr_5_T_1 : _GEN_804; // @[FSM.scala 650:30 FSM.scala 652:27]
  wire [11:0] _GEN_816 = count == 10'h380 ? _L1_rd_addr_6_T_1 : _GEN_805; // @[FSM.scala 650:30 FSM.scala 652:27]
  wire [11:0] _GEN_817 = count == 10'h380 ? _L1_rd_addr_7_T_1 : _GEN_806; // @[FSM.scala 650:30 FSM.scala 652:27]
  wire [11:0] _GEN_818 = count == 10'h380 ? _L1_rd_addr_8_T_1 : _GEN_807; // @[FSM.scala 650:30 FSM.scala 652:27]
  wire [11:0] _GEN_819 = count == 10'h380 ? _L1_rd_addr_9_T_1 : _GEN_808; // @[FSM.scala 650:30 FSM.scala 652:27]
  wire [11:0] _GEN_820 = count == 10'h380 ? _L1_rd_addr_10_T_1 : _GEN_809; // @[FSM.scala 650:30 FSM.scala 652:27]
  wire [11:0] _GEN_821 = count == 10'h380 ? _L1_rd_addr_11_T_1 : _GEN_810; // @[FSM.scala 650:30 FSM.scala 652:27]
  wire  _T_114 = count == 10'h381; // @[FSM.scala 655:20]
  wire [11:0] _GEN_822 = count == 10'h381 ? _L1_rd_addr_2_T_1 : _GEN_812; // @[FSM.scala 655:30 FSM.scala 657:27]
  wire [11:0] _GEN_823 = count == 10'h381 ? _L1_rd_addr_3_T_1 : _GEN_813; // @[FSM.scala 655:30 FSM.scala 657:27]
  wire [11:0] _GEN_824 = count == 10'h381 ? _L1_rd_addr_4_T_1 : _GEN_814; // @[FSM.scala 655:30 FSM.scala 657:27]
  wire [11:0] _GEN_825 = count == 10'h381 ? _L1_rd_addr_5_T_1 : _GEN_815; // @[FSM.scala 655:30 FSM.scala 657:27]
  wire [11:0] _GEN_826 = count == 10'h381 ? _L1_rd_addr_6_T_1 : _GEN_816; // @[FSM.scala 655:30 FSM.scala 657:27]
  wire [11:0] _GEN_827 = count == 10'h381 ? _L1_rd_addr_7_T_1 : _GEN_817; // @[FSM.scala 655:30 FSM.scala 657:27]
  wire [11:0] _GEN_828 = count == 10'h381 ? _L1_rd_addr_8_T_1 : _GEN_818; // @[FSM.scala 655:30 FSM.scala 657:27]
  wire [11:0] _GEN_829 = count == 10'h381 ? _L1_rd_addr_9_T_1 : _GEN_819; // @[FSM.scala 655:30 FSM.scala 657:27]
  wire [11:0] _GEN_830 = count == 10'h381 ? _L1_rd_addr_10_T_1 : _GEN_820; // @[FSM.scala 655:30 FSM.scala 657:27]
  wire [11:0] _GEN_831 = count == 10'h381 ? _L1_rd_addr_11_T_1 : _GEN_821; // @[FSM.scala 655:30 FSM.scala 657:27]
  wire  _T_115 = count == 10'h382; // @[FSM.scala 660:20]
  wire [11:0] _GEN_832 = count == 10'h382 ? _L1_rd_addr_3_T_1 : _GEN_823; // @[FSM.scala 660:30 FSM.scala 662:27]
  wire [11:0] _GEN_833 = count == 10'h382 ? _L1_rd_addr_4_T_1 : _GEN_824; // @[FSM.scala 660:30 FSM.scala 662:27]
  wire [11:0] _GEN_834 = count == 10'h382 ? _L1_rd_addr_5_T_1 : _GEN_825; // @[FSM.scala 660:30 FSM.scala 662:27]
  wire [11:0] _GEN_835 = count == 10'h382 ? _L1_rd_addr_6_T_1 : _GEN_826; // @[FSM.scala 660:30 FSM.scala 662:27]
  wire [11:0] _GEN_836 = count == 10'h382 ? _L1_rd_addr_7_T_1 : _GEN_827; // @[FSM.scala 660:30 FSM.scala 662:27]
  wire [11:0] _GEN_837 = count == 10'h382 ? _L1_rd_addr_8_T_1 : _GEN_828; // @[FSM.scala 660:30 FSM.scala 662:27]
  wire [11:0] _GEN_838 = count == 10'h382 ? _L1_rd_addr_9_T_1 : _GEN_829; // @[FSM.scala 660:30 FSM.scala 662:27]
  wire [11:0] _GEN_839 = count == 10'h382 ? _L1_rd_addr_10_T_1 : _GEN_830; // @[FSM.scala 660:30 FSM.scala 662:27]
  wire [11:0] _GEN_840 = count == 10'h382 ? _L1_rd_addr_11_T_1 : _GEN_831; // @[FSM.scala 660:30 FSM.scala 662:27]
  wire  _T_116 = count == 10'h383; // @[FSM.scala 665:20]
  wire [11:0] _GEN_841 = count == 10'h383 ? _L1_rd_addr_4_T_1 : _GEN_833; // @[FSM.scala 665:30 FSM.scala 667:27]
  wire [11:0] _GEN_842 = count == 10'h383 ? _L1_rd_addr_5_T_1 : _GEN_834; // @[FSM.scala 665:30 FSM.scala 667:27]
  wire [11:0] _GEN_843 = count == 10'h383 ? _L1_rd_addr_6_T_1 : _GEN_835; // @[FSM.scala 665:30 FSM.scala 667:27]
  wire [11:0] _GEN_844 = count == 10'h383 ? _L1_rd_addr_7_T_1 : _GEN_836; // @[FSM.scala 665:30 FSM.scala 667:27]
  wire [11:0] _GEN_845 = count == 10'h383 ? _L1_rd_addr_8_T_1 : _GEN_837; // @[FSM.scala 665:30 FSM.scala 667:27]
  wire [11:0] _GEN_846 = count == 10'h383 ? _L1_rd_addr_9_T_1 : _GEN_838; // @[FSM.scala 665:30 FSM.scala 667:27]
  wire [11:0] _GEN_847 = count == 10'h383 ? _L1_rd_addr_10_T_1 : _GEN_839; // @[FSM.scala 665:30 FSM.scala 667:27]
  wire [11:0] _GEN_848 = count == 10'h383 ? _L1_rd_addr_11_T_1 : _GEN_840; // @[FSM.scala 665:30 FSM.scala 667:27]
  wire  _T_117 = count == 10'h384; // @[FSM.scala 670:20]
  wire [11:0] _GEN_849 = count == 10'h384 ? _L1_rd_addr_5_T_1 : _GEN_842; // @[FSM.scala 670:30 FSM.scala 672:27]
  wire [11:0] _GEN_850 = count == 10'h384 ? _L1_rd_addr_6_T_1 : _GEN_843; // @[FSM.scala 670:30 FSM.scala 672:27]
  wire [11:0] _GEN_851 = count == 10'h384 ? _L1_rd_addr_7_T_1 : _GEN_844; // @[FSM.scala 670:30 FSM.scala 672:27]
  wire [11:0] _GEN_852 = count == 10'h384 ? _L1_rd_addr_8_T_1 : _GEN_845; // @[FSM.scala 670:30 FSM.scala 672:27]
  wire [11:0] _GEN_853 = count == 10'h384 ? _L1_rd_addr_9_T_1 : _GEN_846; // @[FSM.scala 670:30 FSM.scala 672:27]
  wire [11:0] _GEN_854 = count == 10'h384 ? _L1_rd_addr_10_T_1 : _GEN_847; // @[FSM.scala 670:30 FSM.scala 672:27]
  wire [11:0] _GEN_855 = count == 10'h384 ? _L1_rd_addr_11_T_1 : _GEN_848; // @[FSM.scala 670:30 FSM.scala 672:27]
  wire  _T_118 = count == 10'h385; // @[FSM.scala 675:20]
  wire [11:0] _GEN_856 = count == 10'h385 ? _L1_rd_addr_6_T_1 : _GEN_850; // @[FSM.scala 675:30 FSM.scala 677:27]
  wire [11:0] _GEN_857 = count == 10'h385 ? _L1_rd_addr_7_T_1 : _GEN_851; // @[FSM.scala 675:30 FSM.scala 677:27]
  wire [11:0] _GEN_858 = count == 10'h385 ? _L1_rd_addr_8_T_1 : _GEN_852; // @[FSM.scala 675:30 FSM.scala 677:27]
  wire [11:0] _GEN_859 = count == 10'h385 ? _L1_rd_addr_9_T_1 : _GEN_853; // @[FSM.scala 675:30 FSM.scala 677:27]
  wire [11:0] _GEN_860 = count == 10'h385 ? _L1_rd_addr_10_T_1 : _GEN_854; // @[FSM.scala 675:30 FSM.scala 677:27]
  wire [11:0] _GEN_861 = count == 10'h385 ? _L1_rd_addr_11_T_1 : _GEN_855; // @[FSM.scala 675:30 FSM.scala 677:27]
  wire  _T_119 = count == 10'h386; // @[FSM.scala 680:20]
  wire [11:0] _GEN_862 = count == 10'h386 ? _L1_rd_addr_7_T_1 : _GEN_857; // @[FSM.scala 680:30 FSM.scala 682:27]
  wire [11:0] _GEN_863 = count == 10'h386 ? _L1_rd_addr_8_T_1 : _GEN_858; // @[FSM.scala 680:30 FSM.scala 682:27]
  wire [11:0] _GEN_864 = count == 10'h386 ? _L1_rd_addr_9_T_1 : _GEN_859; // @[FSM.scala 680:30 FSM.scala 682:27]
  wire [11:0] _GEN_865 = count == 10'h386 ? _L1_rd_addr_10_T_1 : _GEN_860; // @[FSM.scala 680:30 FSM.scala 682:27]
  wire [11:0] _GEN_866 = count == 10'h386 ? _L1_rd_addr_11_T_1 : _GEN_861; // @[FSM.scala 680:30 FSM.scala 682:27]
  wire  _T_120 = count == 10'h387; // @[FSM.scala 685:20]
  wire [11:0] _GEN_867 = count == 10'h387 ? _L1_rd_addr_8_T_1 : _GEN_863; // @[FSM.scala 685:30 FSM.scala 687:27]
  wire [11:0] _GEN_868 = count == 10'h387 ? _L1_rd_addr_9_T_1 : _GEN_864; // @[FSM.scala 685:30 FSM.scala 687:27]
  wire [11:0] _GEN_869 = count == 10'h387 ? _L1_rd_addr_10_T_1 : _GEN_865; // @[FSM.scala 685:30 FSM.scala 687:27]
  wire [11:0] _GEN_870 = count == 10'h387 ? _L1_rd_addr_11_T_1 : _GEN_866; // @[FSM.scala 685:30 FSM.scala 687:27]
  wire  _T_121 = count == 10'h388; // @[FSM.scala 690:20]
  wire [11:0] _GEN_871 = count == 10'h388 ? _L1_rd_addr_9_T_1 : _GEN_868; // @[FSM.scala 690:30 FSM.scala 692:27]
  wire [11:0] _GEN_872 = count == 10'h388 ? _L1_rd_addr_10_T_1 : _GEN_869; // @[FSM.scala 690:30 FSM.scala 692:27]
  wire [11:0] _GEN_873 = count == 10'h388 ? _L1_rd_addr_11_T_1 : _GEN_870; // @[FSM.scala 690:30 FSM.scala 692:27]
  wire  _T_122 = count == 10'h389; // @[FSM.scala 695:20]
  wire [11:0] _GEN_874 = count == 10'h389 ? _L1_rd_addr_10_T_1 : _GEN_872; // @[FSM.scala 695:30 FSM.scala 697:27]
  wire [11:0] _GEN_875 = count == 10'h389 ? _L1_rd_addr_11_T_1 : _GEN_873; // @[FSM.scala 695:30 FSM.scala 697:27]
  wire  _T_123 = count == 10'h38a; // @[FSM.scala 700:20]
  wire [11:0] _GEN_876 = count == 10'h38a ? _L1_rd_addr_11_T_1 : _GEN_875; // @[FSM.scala 700:30 FSM.scala 702:27]
  wire  _T_124 = count >= 10'he; // @[FSM.scala 706:21]
  wire  _T_126 = count >= 10'he & count <= 10'h38d; // @[FSM.scala 706:30]
  wire  _T_127 = count1 == 7'he; // @[FSM.scala 707:23]
  wire [5:0] _Zt_wrAddr_T_1 = Zt_wrAddr + 6'h1; // @[FSM.scala 712:36]
  wire [5:0] _GEN_877 = count1 == 7'he ? 6'h0 : _Zt_wrAddr_T_1; // @[FSM.scala 707:33 FSM.scala 708:23 FSM.scala 712:23]
  wire [5:0] _GEN_879 = count >= 10'he & count <= 10'h38d ? _GEN_877 : _GEN_722; // @[FSM.scala 706:50]
  wire  _GEN_880 = count >= 10'he & count <= 10'h38d | Zt_wrEna; // @[FSM.scala 706:50 FSM.scala 82:36]
  wire  _T_128 = count == 10'h38e; // @[FSM.scala 717:20]
  wire [9:0] _GEN_881 = count == 10'h38e ? 10'h0 : _GEN_701; // @[FSM.scala 717:30 FSM.scala 718:17]
  wire [6:0] _GEN_882 = count == 10'h38e ? 7'h0 : _GEN_702; // @[FSM.scala 717:30 FSM.scala 719:18]
  wire  _GEN_883 = count == 10'h38e ? 1'h0 : _GEN_880; // @[FSM.scala 717:30 FSM.scala 720:20]
  wire [3:0] _GEN_884 = count == 10'h38e ? 4'h2 : _GEN_700; // @[FSM.scala 717:30 FSM.scala 721:21]
  wire [9:0] _GEN_885 = gru_state == 4'h1 ? _GEN_881 : _GEN_678; // @[FSM.scala 543:30]
  wire [6:0] _GEN_886 = gru_state == 4'h1 ? _GEN_882 : count1; // @[FSM.scala 543:30 FSM.scala 162:23]
  wire [2:0] _GEN_887 = gru_state == 4'h1 ? _GEN_725 : _GEN_679; // @[FSM.scala 543:30]
  wire [9:0] _GEN_888 = gru_state == 4'h1 ? _GEN_726 : _GEN_681; // @[FSM.scala 543:30]
  wire [5:0] _GEN_889 = gru_state == 4'h1 ? _GEN_727 : _GEN_682; // @[FSM.scala 543:30]
  wire [11:0] _GEN_890 = gru_state == 4'h1 ? _GEN_732 : _GEN_680; // @[FSM.scala 543:30]
  wire [7:0] _GEN_891 = gru_state == 4'h1 ? _GEN_729 : PEArray_ctrl_2_gru_out_width; // @[FSM.scala 543:30 FSM.scala 64:28]
  wire [11:0] _GEN_892 = gru_state == 4'h1 ? _GEN_799 : _GEN_688; // @[FSM.scala 543:30]
  wire [11:0] _GEN_893 = gru_state == 4'h1 ? _GEN_811 : _GEN_689; // @[FSM.scala 543:30]
  wire [11:0] _GEN_894 = gru_state == 4'h1 ? _GEN_822 : _GEN_690; // @[FSM.scala 543:30]
  wire [11:0] _GEN_895 = gru_state == 4'h1 ? _GEN_832 : _GEN_691; // @[FSM.scala 543:30]
  wire [11:0] _GEN_896 = gru_state == 4'h1 ? _GEN_841 : _GEN_692; // @[FSM.scala 543:30]
  wire [11:0] _GEN_897 = gru_state == 4'h1 ? _GEN_849 : _GEN_693; // @[FSM.scala 543:30]
  wire [11:0] _GEN_898 = gru_state == 4'h1 ? _GEN_856 : _GEN_694; // @[FSM.scala 543:30]
  wire [11:0] _GEN_899 = gru_state == 4'h1 ? _GEN_862 : _GEN_695; // @[FSM.scala 543:30]
  wire [11:0] _GEN_900 = gru_state == 4'h1 ? _GEN_867 : _GEN_696; // @[FSM.scala 543:30]
  wire [11:0] _GEN_901 = gru_state == 4'h1 ? _GEN_871 : _GEN_697; // @[FSM.scala 543:30]
  wire [11:0] _GEN_902 = gru_state == 4'h1 ? _GEN_874 : _GEN_698; // @[FSM.scala 543:30]
  wire [11:0] _GEN_903 = gru_state == 4'h1 ? _GEN_876 : _GEN_699; // @[FSM.scala 543:30]
  wire [1:0] _GEN_904 = gru_state == 4'h1 ? _GEN_720 : _GEN_683; // @[FSM.scala 543:30]
  wire [3:0] _GEN_905 = gru_state == 4'h1 ? _GEN_721 : _GEN_684; // @[FSM.scala 543:30]
  wire [5:0] _GEN_906 = gru_state == 4'h1 ? _GEN_879 : Zt_wrAddr; // @[FSM.scala 543:30 FSM.scala 83:36]
  wire [1:0] _GEN_907 = gru_state == 4'h1 ? _GEN_723 : BN_Unit_ctrl; // @[FSM.scala 543:30 FSM.scala 69:28]
  wire [1:0] _GEN_908 = gru_state == 4'h1 ? _GEN_724 : Activation_ctrl; // @[FSM.scala 543:30 FSM.scala 75:32]
  wire [11:0] _GEN_909 = gru_state == 4'h1 ? _GEN_730 : _GEN_685; // @[FSM.scala 543:30]
  wire [11:0] _GEN_910 = gru_state == 4'h1 ? _GEN_731 : _GEN_686; // @[FSM.scala 543:30]
  wire  _GEN_911 = gru_state == 4'h1 ? _GEN_883 : Zt_wrEna; // @[FSM.scala 543:30 FSM.scala 82:36]
  wire [3:0] _GEN_912 = gru_state == 4'h1 ? _GEN_884 : _GEN_700; // @[FSM.scala 543:30]
  wire [9:0] _GEN_913 = _T_92 ? _count_T_1 : _GEN_885; // @[FSM.scala 726:30 FSM.scala 727:17]
  wire [2:0] _GEN_915 = _T_3 ? 3'h4 : _GEN_887; // @[FSM.scala 736:28 FSM.scala 738:35]
  wire [9:0] _GEN_916 = _T_3 ? 10'h37f : _GEN_888; // @[FSM.scala 736:28 FSM.scala 739:33]
  wire [5:0] _GEN_917 = _T_3 ? 6'hf : _GEN_889; // @[FSM.scala 736:28 FSM.scala 740:35]
  wire [11:0] _GEN_918 = _T_3 ? 12'h800 : _GEN_890; // @[FSM.scala 736:28 FSM.scala 741:32]
  wire [7:0] _GEN_919 = _T_3 ? 8'h40 : _GEN_891; // @[FSM.scala 736:28 FSM.scala 742:41]
  wire [1:0] _GEN_920 = _T_3 ? 2'h0 : _GEN_904; // @[FSM.scala 736:28 FSM.scala 745:30]
  wire [3:0] _GEN_921 = _T_3 ? 4'h0 : _GEN_905; // @[FSM.scala 736:28 FSM.scala 746:26]
  wire [5:0] _GEN_922 = _T_3 ? 6'h0 : Rt_wrAddr; // @[FSM.scala 736:28 FSM.scala 749:21 FSM.scala 86:36]
  wire [1:0] _GEN_923 = _T_3 ? 2'h2 : _GEN_907; // @[FSM.scala 736:28 FSM.scala 750:24]
  wire [1:0] _GEN_924 = _T_3 ? 2'h1 : _GEN_908; // @[FSM.scala 736:28 FSM.scala 751:27]
  wire [2:0] _GEN_925 = _T_39 ? 3'h4 : _GEN_915; // @[FSM.scala 755:48 FSM.scala 756:35]
  wire [9:0] _GEN_926 = _T_39 ? 10'h37f : _GEN_916; // @[FSM.scala 755:48 FSM.scala 757:33]
  wire [5:0] _GEN_927 = _T_39 ? 6'hf : _GEN_917; // @[FSM.scala 755:48 FSM.scala 758:35]
  wire [11:0] _GEN_928 = _T_39 ? {{1'd0}, PEArray_ctrl_2_mask[11:1]} : _GEN_918; // @[FSM.scala 755:48 FSM.scala 759:32]
  wire [7:0] _GEN_929 = _T_39 ? 8'h40 : _GEN_919; // @[FSM.scala 755:48 FSM.scala 760:41]
  wire [11:0] _GEN_930 = _T_40 ? 12'h0 : _GEN_909; // @[FSM.scala 762:29 FSM.scala 764:34]
  wire [11:0] _GEN_931 = _T_40 ? 12'h0 : _GEN_910; // @[FSM.scala 762:29 FSM.scala 764:34]
  wire [11:0] _GEN_932 = _T_40 ? 12'h0 : _GEN_928; // @[FSM.scala 762:29 FSM.scala 764:34]
  wire [11:0] _GEN_933 = _T_5 ? _L1_rd_addr_0_T_1 : _GEN_892; // @[FSM.scala 769:28 FSM.scala 771:27]
  wire [11:0] _GEN_934 = _T_48 ? _L1_rd_addr_0_T_1 : _GEN_933; // @[FSM.scala 774:28 FSM.scala 776:27]
  wire [11:0] _GEN_935 = _T_48 ? _L1_rd_addr_1_T_1 : _GEN_893; // @[FSM.scala 774:28 FSM.scala 776:27]
  wire [11:0] _GEN_936 = _T_49 ? _L1_rd_addr_0_T_1 : _GEN_934; // @[FSM.scala 779:28 FSM.scala 781:27]
  wire [11:0] _GEN_937 = _T_49 ? _L1_rd_addr_1_T_1 : _GEN_935; // @[FSM.scala 779:28 FSM.scala 781:27]
  wire [11:0] _GEN_938 = _T_49 ? _L1_rd_addr_2_T_1 : _GEN_894; // @[FSM.scala 779:28 FSM.scala 781:27]
  wire [11:0] _GEN_939 = _T_21 ? _L1_rd_addr_0_T_1 : _GEN_936; // @[FSM.scala 784:28 FSM.scala 786:27]
  wire [11:0] _GEN_940 = _T_21 ? _L1_rd_addr_1_T_1 : _GEN_937; // @[FSM.scala 784:28 FSM.scala 786:27]
  wire [11:0] _GEN_941 = _T_21 ? _L1_rd_addr_2_T_1 : _GEN_938; // @[FSM.scala 784:28 FSM.scala 786:27]
  wire [11:0] _GEN_942 = _T_21 ? _L1_rd_addr_3_T_1 : _GEN_895; // @[FSM.scala 784:28 FSM.scala 786:27]
  wire [11:0] _GEN_943 = _T_51 ? _L1_rd_addr_0_T_1 : _GEN_939; // @[FSM.scala 789:28 FSM.scala 791:27]
  wire [11:0] _GEN_944 = _T_51 ? _L1_rd_addr_1_T_1 : _GEN_940; // @[FSM.scala 789:28 FSM.scala 791:27]
  wire [11:0] _GEN_945 = _T_51 ? _L1_rd_addr_2_T_1 : _GEN_941; // @[FSM.scala 789:28 FSM.scala 791:27]
  wire [11:0] _GEN_946 = _T_51 ? _L1_rd_addr_3_T_1 : _GEN_942; // @[FSM.scala 789:28 FSM.scala 791:27]
  wire [11:0] _GEN_947 = _T_51 ? _L1_rd_addr_4_T_1 : _GEN_896; // @[FSM.scala 789:28 FSM.scala 791:27]
  wire [11:0] _GEN_948 = _T_52 ? _L1_rd_addr_0_T_1 : _GEN_943; // @[FSM.scala 794:28 FSM.scala 796:27]
  wire [11:0] _GEN_949 = _T_52 ? _L1_rd_addr_1_T_1 : _GEN_944; // @[FSM.scala 794:28 FSM.scala 796:27]
  wire [11:0] _GEN_950 = _T_52 ? _L1_rd_addr_2_T_1 : _GEN_945; // @[FSM.scala 794:28 FSM.scala 796:27]
  wire [11:0] _GEN_951 = _T_52 ? _L1_rd_addr_3_T_1 : _GEN_946; // @[FSM.scala 794:28 FSM.scala 796:27]
  wire [11:0] _GEN_952 = _T_52 ? _L1_rd_addr_4_T_1 : _GEN_947; // @[FSM.scala 794:28 FSM.scala 796:27]
  wire [11:0] _GEN_953 = _T_52 ? _L1_rd_addr_5_T_1 : _GEN_897; // @[FSM.scala 794:28 FSM.scala 796:27]
  wire [11:0] _GEN_954 = _T_53 ? _L1_rd_addr_0_T_1 : _GEN_948; // @[FSM.scala 799:28 FSM.scala 801:27]
  wire [11:0] _GEN_955 = _T_53 ? _L1_rd_addr_1_T_1 : _GEN_949; // @[FSM.scala 799:28 FSM.scala 801:27]
  wire [11:0] _GEN_956 = _T_53 ? _L1_rd_addr_2_T_1 : _GEN_950; // @[FSM.scala 799:28 FSM.scala 801:27]
  wire [11:0] _GEN_957 = _T_53 ? _L1_rd_addr_3_T_1 : _GEN_951; // @[FSM.scala 799:28 FSM.scala 801:27]
  wire [11:0] _GEN_958 = _T_53 ? _L1_rd_addr_4_T_1 : _GEN_952; // @[FSM.scala 799:28 FSM.scala 801:27]
  wire [11:0] _GEN_959 = _T_53 ? _L1_rd_addr_5_T_1 : _GEN_953; // @[FSM.scala 799:28 FSM.scala 801:27]
  wire [11:0] _GEN_960 = _T_53 ? _L1_rd_addr_6_T_1 : _GEN_898; // @[FSM.scala 799:28 FSM.scala 801:27]
  wire [11:0] _GEN_961 = _T_54 ? _L1_rd_addr_0_T_1 : _GEN_954; // @[FSM.scala 804:28 FSM.scala 806:27]
  wire [11:0] _GEN_962 = _T_54 ? _L1_rd_addr_1_T_1 : _GEN_955; // @[FSM.scala 804:28 FSM.scala 806:27]
  wire [11:0] _GEN_963 = _T_54 ? _L1_rd_addr_2_T_1 : _GEN_956; // @[FSM.scala 804:28 FSM.scala 806:27]
  wire [11:0] _GEN_964 = _T_54 ? _L1_rd_addr_3_T_1 : _GEN_957; // @[FSM.scala 804:28 FSM.scala 806:27]
  wire [11:0] _GEN_965 = _T_54 ? _L1_rd_addr_4_T_1 : _GEN_958; // @[FSM.scala 804:28 FSM.scala 806:27]
  wire [11:0] _GEN_966 = _T_54 ? _L1_rd_addr_5_T_1 : _GEN_959; // @[FSM.scala 804:28 FSM.scala 806:27]
  wire [11:0] _GEN_967 = _T_54 ? _L1_rd_addr_6_T_1 : _GEN_960; // @[FSM.scala 804:28 FSM.scala 806:27]
  wire [11:0] _GEN_968 = _T_54 ? _L1_rd_addr_7_T_1 : _GEN_899; // @[FSM.scala 804:28 FSM.scala 806:27]
  wire [11:0] _GEN_969 = _T_55 ? _L1_rd_addr_0_T_1 : _GEN_961; // @[FSM.scala 809:28 FSM.scala 811:27]
  wire [11:0] _GEN_970 = _T_55 ? _L1_rd_addr_1_T_1 : _GEN_962; // @[FSM.scala 809:28 FSM.scala 811:27]
  wire [11:0] _GEN_971 = _T_55 ? _L1_rd_addr_2_T_1 : _GEN_963; // @[FSM.scala 809:28 FSM.scala 811:27]
  wire [11:0] _GEN_972 = _T_55 ? _L1_rd_addr_3_T_1 : _GEN_964; // @[FSM.scala 809:28 FSM.scala 811:27]
  wire [11:0] _GEN_973 = _T_55 ? _L1_rd_addr_4_T_1 : _GEN_965; // @[FSM.scala 809:28 FSM.scala 811:27]
  wire [11:0] _GEN_974 = _T_55 ? _L1_rd_addr_5_T_1 : _GEN_966; // @[FSM.scala 809:28 FSM.scala 811:27]
  wire [11:0] _GEN_975 = _T_55 ? _L1_rd_addr_6_T_1 : _GEN_967; // @[FSM.scala 809:28 FSM.scala 811:27]
  wire [11:0] _GEN_976 = _T_55 ? _L1_rd_addr_7_T_1 : _GEN_968; // @[FSM.scala 809:28 FSM.scala 811:27]
  wire [11:0] _GEN_977 = _T_55 ? _L1_rd_addr_8_T_1 : _GEN_900; // @[FSM.scala 809:28 FSM.scala 811:27]
  wire [11:0] _GEN_978 = _T_56 ? _L1_rd_addr_0_T_1 : _GEN_969; // @[FSM.scala 814:29 FSM.scala 816:27]
  wire [11:0] _GEN_979 = _T_56 ? _L1_rd_addr_1_T_1 : _GEN_970; // @[FSM.scala 814:29 FSM.scala 816:27]
  wire [11:0] _GEN_980 = _T_56 ? _L1_rd_addr_2_T_1 : _GEN_971; // @[FSM.scala 814:29 FSM.scala 816:27]
  wire [11:0] _GEN_981 = _T_56 ? _L1_rd_addr_3_T_1 : _GEN_972; // @[FSM.scala 814:29 FSM.scala 816:27]
  wire [11:0] _GEN_982 = _T_56 ? _L1_rd_addr_4_T_1 : _GEN_973; // @[FSM.scala 814:29 FSM.scala 816:27]
  wire [11:0] _GEN_983 = _T_56 ? _L1_rd_addr_5_T_1 : _GEN_974; // @[FSM.scala 814:29 FSM.scala 816:27]
  wire [11:0] _GEN_984 = _T_56 ? _L1_rd_addr_6_T_1 : _GEN_975; // @[FSM.scala 814:29 FSM.scala 816:27]
  wire [11:0] _GEN_985 = _T_56 ? _L1_rd_addr_7_T_1 : _GEN_976; // @[FSM.scala 814:29 FSM.scala 816:27]
  wire [11:0] _GEN_986 = _T_56 ? _L1_rd_addr_8_T_1 : _GEN_977; // @[FSM.scala 814:29 FSM.scala 816:27]
  wire [11:0] _GEN_987 = _T_56 ? _L1_rd_addr_9_T_1 : _GEN_901; // @[FSM.scala 814:29 FSM.scala 816:27]
  wire [11:0] _GEN_988 = _T_57 ? _L1_rd_addr_0_T_1 : _GEN_978; // @[FSM.scala 819:29 FSM.scala 821:27]
  wire [11:0] _GEN_989 = _T_57 ? _L1_rd_addr_1_T_1 : _GEN_979; // @[FSM.scala 819:29 FSM.scala 821:27]
  wire [11:0] _GEN_990 = _T_57 ? _L1_rd_addr_2_T_1 : _GEN_980; // @[FSM.scala 819:29 FSM.scala 821:27]
  wire [11:0] _GEN_991 = _T_57 ? _L1_rd_addr_3_T_1 : _GEN_981; // @[FSM.scala 819:29 FSM.scala 821:27]
  wire [11:0] _GEN_992 = _T_57 ? _L1_rd_addr_4_T_1 : _GEN_982; // @[FSM.scala 819:29 FSM.scala 821:27]
  wire [11:0] _GEN_993 = _T_57 ? _L1_rd_addr_5_T_1 : _GEN_983; // @[FSM.scala 819:29 FSM.scala 821:27]
  wire [11:0] _GEN_994 = _T_57 ? _L1_rd_addr_6_T_1 : _GEN_984; // @[FSM.scala 819:29 FSM.scala 821:27]
  wire [11:0] _GEN_995 = _T_57 ? _L1_rd_addr_7_T_1 : _GEN_985; // @[FSM.scala 819:29 FSM.scala 821:27]
  wire [11:0] _GEN_996 = _T_57 ? _L1_rd_addr_8_T_1 : _GEN_986; // @[FSM.scala 819:29 FSM.scala 821:27]
  wire [11:0] _GEN_997 = _T_57 ? _L1_rd_addr_9_T_1 : _GEN_987; // @[FSM.scala 819:29 FSM.scala 821:27]
  wire [11:0] _GEN_998 = _T_57 ? _L1_rd_addr_10_T_1 : _GEN_902; // @[FSM.scala 819:29 FSM.scala 821:27]
  wire [11:0] _GEN_999 = _T_112 ? _L1_rd_addr_0_T_1 : _GEN_988; // @[FSM.scala 824:50 FSM.scala 826:27]
  wire [11:0] _GEN_1000 = _T_112 ? _L1_rd_addr_1_T_1 : _GEN_989; // @[FSM.scala 824:50 FSM.scala 826:27]
  wire [11:0] _GEN_1001 = _T_112 ? _L1_rd_addr_2_T_1 : _GEN_990; // @[FSM.scala 824:50 FSM.scala 826:27]
  wire [11:0] _GEN_1002 = _T_112 ? _L1_rd_addr_3_T_1 : _GEN_991; // @[FSM.scala 824:50 FSM.scala 826:27]
  wire [11:0] _GEN_1003 = _T_112 ? _L1_rd_addr_4_T_1 : _GEN_992; // @[FSM.scala 824:50 FSM.scala 826:27]
  wire [11:0] _GEN_1004 = _T_112 ? _L1_rd_addr_5_T_1 : _GEN_993; // @[FSM.scala 824:50 FSM.scala 826:27]
  wire [11:0] _GEN_1005 = _T_112 ? _L1_rd_addr_6_T_1 : _GEN_994; // @[FSM.scala 824:50 FSM.scala 826:27]
  wire [11:0] _GEN_1006 = _T_112 ? _L1_rd_addr_7_T_1 : _GEN_995; // @[FSM.scala 824:50 FSM.scala 826:27]
  wire [11:0] _GEN_1007 = _T_112 ? _L1_rd_addr_8_T_1 : _GEN_996; // @[FSM.scala 824:50 FSM.scala 826:27]
  wire [11:0] _GEN_1008 = _T_112 ? _L1_rd_addr_9_T_1 : _GEN_997; // @[FSM.scala 824:50 FSM.scala 826:27]
  wire [11:0] _GEN_1009 = _T_112 ? _L1_rd_addr_10_T_1 : _GEN_998; // @[FSM.scala 824:50 FSM.scala 826:27]
  wire [11:0] _GEN_1010 = _T_112 ? _L1_rd_addr_11_T_1 : _GEN_903; // @[FSM.scala 824:50 FSM.scala 826:27]
  wire [11:0] _GEN_1011 = _T_113 ? _L1_rd_addr_1_T_1 : _GEN_1000; // @[FSM.scala 829:30 FSM.scala 831:27]
  wire [11:0] _GEN_1012 = _T_113 ? _L1_rd_addr_2_T_1 : _GEN_1001; // @[FSM.scala 829:30 FSM.scala 831:27]
  wire [11:0] _GEN_1013 = _T_113 ? _L1_rd_addr_3_T_1 : _GEN_1002; // @[FSM.scala 829:30 FSM.scala 831:27]
  wire [11:0] _GEN_1014 = _T_113 ? _L1_rd_addr_4_T_1 : _GEN_1003; // @[FSM.scala 829:30 FSM.scala 831:27]
  wire [11:0] _GEN_1015 = _T_113 ? _L1_rd_addr_5_T_1 : _GEN_1004; // @[FSM.scala 829:30 FSM.scala 831:27]
  wire [11:0] _GEN_1016 = _T_113 ? _L1_rd_addr_6_T_1 : _GEN_1005; // @[FSM.scala 829:30 FSM.scala 831:27]
  wire [11:0] _GEN_1017 = _T_113 ? _L1_rd_addr_7_T_1 : _GEN_1006; // @[FSM.scala 829:30 FSM.scala 831:27]
  wire [11:0] _GEN_1018 = _T_113 ? _L1_rd_addr_8_T_1 : _GEN_1007; // @[FSM.scala 829:30 FSM.scala 831:27]
  wire [11:0] _GEN_1019 = _T_113 ? _L1_rd_addr_9_T_1 : _GEN_1008; // @[FSM.scala 829:30 FSM.scala 831:27]
  wire [11:0] _GEN_1020 = _T_113 ? _L1_rd_addr_10_T_1 : _GEN_1009; // @[FSM.scala 829:30 FSM.scala 831:27]
  wire [11:0] _GEN_1021 = _T_113 ? _L1_rd_addr_11_T_1 : _GEN_1010; // @[FSM.scala 829:30 FSM.scala 831:27]
  wire [11:0] _GEN_1022 = _T_114 ? _L1_rd_addr_2_T_1 : _GEN_1012; // @[FSM.scala 834:30 FSM.scala 836:27]
  wire [11:0] _GEN_1023 = _T_114 ? _L1_rd_addr_3_T_1 : _GEN_1013; // @[FSM.scala 834:30 FSM.scala 836:27]
  wire [11:0] _GEN_1024 = _T_114 ? _L1_rd_addr_4_T_1 : _GEN_1014; // @[FSM.scala 834:30 FSM.scala 836:27]
  wire [11:0] _GEN_1025 = _T_114 ? _L1_rd_addr_5_T_1 : _GEN_1015; // @[FSM.scala 834:30 FSM.scala 836:27]
  wire [11:0] _GEN_1026 = _T_114 ? _L1_rd_addr_6_T_1 : _GEN_1016; // @[FSM.scala 834:30 FSM.scala 836:27]
  wire [11:0] _GEN_1027 = _T_114 ? _L1_rd_addr_7_T_1 : _GEN_1017; // @[FSM.scala 834:30 FSM.scala 836:27]
  wire [11:0] _GEN_1028 = _T_114 ? _L1_rd_addr_8_T_1 : _GEN_1018; // @[FSM.scala 834:30 FSM.scala 836:27]
  wire [11:0] _GEN_1029 = _T_114 ? _L1_rd_addr_9_T_1 : _GEN_1019; // @[FSM.scala 834:30 FSM.scala 836:27]
  wire [11:0] _GEN_1030 = _T_114 ? _L1_rd_addr_10_T_1 : _GEN_1020; // @[FSM.scala 834:30 FSM.scala 836:27]
  wire [11:0] _GEN_1031 = _T_114 ? _L1_rd_addr_11_T_1 : _GEN_1021; // @[FSM.scala 834:30 FSM.scala 836:27]
  wire [11:0] _GEN_1032 = _T_115 ? _L1_rd_addr_3_T_1 : _GEN_1023; // @[FSM.scala 839:30 FSM.scala 841:27]
  wire [11:0] _GEN_1033 = _T_115 ? _L1_rd_addr_4_T_1 : _GEN_1024; // @[FSM.scala 839:30 FSM.scala 841:27]
  wire [11:0] _GEN_1034 = _T_115 ? _L1_rd_addr_5_T_1 : _GEN_1025; // @[FSM.scala 839:30 FSM.scala 841:27]
  wire [11:0] _GEN_1035 = _T_115 ? _L1_rd_addr_6_T_1 : _GEN_1026; // @[FSM.scala 839:30 FSM.scala 841:27]
  wire [11:0] _GEN_1036 = _T_115 ? _L1_rd_addr_7_T_1 : _GEN_1027; // @[FSM.scala 839:30 FSM.scala 841:27]
  wire [11:0] _GEN_1037 = _T_115 ? _L1_rd_addr_8_T_1 : _GEN_1028; // @[FSM.scala 839:30 FSM.scala 841:27]
  wire [11:0] _GEN_1038 = _T_115 ? _L1_rd_addr_9_T_1 : _GEN_1029; // @[FSM.scala 839:30 FSM.scala 841:27]
  wire [11:0] _GEN_1039 = _T_115 ? _L1_rd_addr_10_T_1 : _GEN_1030; // @[FSM.scala 839:30 FSM.scala 841:27]
  wire [11:0] _GEN_1040 = _T_115 ? _L1_rd_addr_11_T_1 : _GEN_1031; // @[FSM.scala 839:30 FSM.scala 841:27]
  wire [11:0] _GEN_1041 = _T_116 ? _L1_rd_addr_4_T_1 : _GEN_1033; // @[FSM.scala 844:30 FSM.scala 846:27]
  wire [11:0] _GEN_1042 = _T_116 ? _L1_rd_addr_5_T_1 : _GEN_1034; // @[FSM.scala 844:30 FSM.scala 846:27]
  wire [11:0] _GEN_1043 = _T_116 ? _L1_rd_addr_6_T_1 : _GEN_1035; // @[FSM.scala 844:30 FSM.scala 846:27]
  wire [11:0] _GEN_1044 = _T_116 ? _L1_rd_addr_7_T_1 : _GEN_1036; // @[FSM.scala 844:30 FSM.scala 846:27]
  wire [11:0] _GEN_1045 = _T_116 ? _L1_rd_addr_8_T_1 : _GEN_1037; // @[FSM.scala 844:30 FSM.scala 846:27]
  wire [11:0] _GEN_1046 = _T_116 ? _L1_rd_addr_9_T_1 : _GEN_1038; // @[FSM.scala 844:30 FSM.scala 846:27]
  wire [11:0] _GEN_1047 = _T_116 ? _L1_rd_addr_10_T_1 : _GEN_1039; // @[FSM.scala 844:30 FSM.scala 846:27]
  wire [11:0] _GEN_1048 = _T_116 ? _L1_rd_addr_11_T_1 : _GEN_1040; // @[FSM.scala 844:30 FSM.scala 846:27]
  wire [11:0] _GEN_1049 = _T_117 ? _L1_rd_addr_5_T_1 : _GEN_1042; // @[FSM.scala 849:30 FSM.scala 851:27]
  wire [11:0] _GEN_1050 = _T_117 ? _L1_rd_addr_6_T_1 : _GEN_1043; // @[FSM.scala 849:30 FSM.scala 851:27]
  wire [11:0] _GEN_1051 = _T_117 ? _L1_rd_addr_7_T_1 : _GEN_1044; // @[FSM.scala 849:30 FSM.scala 851:27]
  wire [11:0] _GEN_1052 = _T_117 ? _L1_rd_addr_8_T_1 : _GEN_1045; // @[FSM.scala 849:30 FSM.scala 851:27]
  wire [11:0] _GEN_1053 = _T_117 ? _L1_rd_addr_9_T_1 : _GEN_1046; // @[FSM.scala 849:30 FSM.scala 851:27]
  wire [11:0] _GEN_1054 = _T_117 ? _L1_rd_addr_10_T_1 : _GEN_1047; // @[FSM.scala 849:30 FSM.scala 851:27]
  wire [11:0] _GEN_1055 = _T_117 ? _L1_rd_addr_11_T_1 : _GEN_1048; // @[FSM.scala 849:30 FSM.scala 851:27]
  wire [11:0] _GEN_1056 = _T_118 ? _L1_rd_addr_6_T_1 : _GEN_1050; // @[FSM.scala 854:30 FSM.scala 856:27]
  wire [11:0] _GEN_1057 = _T_118 ? _L1_rd_addr_7_T_1 : _GEN_1051; // @[FSM.scala 854:30 FSM.scala 856:27]
  wire [11:0] _GEN_1058 = _T_118 ? _L1_rd_addr_8_T_1 : _GEN_1052; // @[FSM.scala 854:30 FSM.scala 856:27]
  wire [11:0] _GEN_1059 = _T_118 ? _L1_rd_addr_9_T_1 : _GEN_1053; // @[FSM.scala 854:30 FSM.scala 856:27]
  wire [11:0] _GEN_1060 = _T_118 ? _L1_rd_addr_10_T_1 : _GEN_1054; // @[FSM.scala 854:30 FSM.scala 856:27]
  wire [11:0] _GEN_1061 = _T_118 ? _L1_rd_addr_11_T_1 : _GEN_1055; // @[FSM.scala 854:30 FSM.scala 856:27]
  wire [11:0] _GEN_1062 = _T_119 ? _L1_rd_addr_7_T_1 : _GEN_1057; // @[FSM.scala 859:30 FSM.scala 861:27]
  wire [11:0] _GEN_1063 = _T_119 ? _L1_rd_addr_8_T_1 : _GEN_1058; // @[FSM.scala 859:30 FSM.scala 861:27]
  wire [11:0] _GEN_1064 = _T_119 ? _L1_rd_addr_9_T_1 : _GEN_1059; // @[FSM.scala 859:30 FSM.scala 861:27]
  wire [11:0] _GEN_1065 = _T_119 ? _L1_rd_addr_10_T_1 : _GEN_1060; // @[FSM.scala 859:30 FSM.scala 861:27]
  wire [11:0] _GEN_1066 = _T_119 ? _L1_rd_addr_11_T_1 : _GEN_1061; // @[FSM.scala 859:30 FSM.scala 861:27]
  wire [11:0] _GEN_1067 = _T_120 ? _L1_rd_addr_8_T_1 : _GEN_1063; // @[FSM.scala 864:30 FSM.scala 866:27]
  wire [11:0] _GEN_1068 = _T_120 ? _L1_rd_addr_9_T_1 : _GEN_1064; // @[FSM.scala 864:30 FSM.scala 866:27]
  wire [11:0] _GEN_1069 = _T_120 ? _L1_rd_addr_10_T_1 : _GEN_1065; // @[FSM.scala 864:30 FSM.scala 866:27]
  wire [11:0] _GEN_1070 = _T_120 ? _L1_rd_addr_11_T_1 : _GEN_1066; // @[FSM.scala 864:30 FSM.scala 866:27]
  wire [11:0] _GEN_1071 = _T_121 ? _L1_rd_addr_9_T_1 : _GEN_1068; // @[FSM.scala 869:30 FSM.scala 871:27]
  wire [11:0] _GEN_1072 = _T_121 ? _L1_rd_addr_10_T_1 : _GEN_1069; // @[FSM.scala 869:30 FSM.scala 871:27]
  wire [11:0] _GEN_1073 = _T_121 ? _L1_rd_addr_11_T_1 : _GEN_1070; // @[FSM.scala 869:30 FSM.scala 871:27]
  wire [11:0] _GEN_1074 = _T_122 ? _L1_rd_addr_10_T_1 : _GEN_1072; // @[FSM.scala 874:30 FSM.scala 876:27]
  wire [11:0] _GEN_1075 = _T_122 ? _L1_rd_addr_11_T_1 : _GEN_1073; // @[FSM.scala 874:30 FSM.scala 876:27]
  wire [11:0] _GEN_1076 = _T_123 ? _L1_rd_addr_11_T_1 : _GEN_1075; // @[FSM.scala 879:30 FSM.scala 881:27]
  wire [5:0] _Rt_wrAddr_T_1 = Rt_wrAddr + 6'h1; // @[FSM.scala 891:38]
  wire [5:0] _GEN_1077 = _T_127 ? 6'h0 : _Rt_wrAddr_T_1; // @[FSM.scala 886:33 FSM.scala 887:23 FSM.scala 891:25]
  wire [5:0] _GEN_1079 = _T_126 ? _GEN_1077 : _GEN_922; // @[FSM.scala 885:50]
  wire  _GEN_1080 = _T_126 | Rt_wrEna; // @[FSM.scala 885:50 FSM.scala 85:36]
  wire [9:0] _GEN_1081 = _T_128 ? 10'h0 : _GEN_913; // @[FSM.scala 896:30 FSM.scala 897:17]
  wire  _GEN_1083 = _T_128 ? 1'h0 : _GEN_1080; // @[FSM.scala 896:30 FSM.scala 899:20]
  wire [3:0] _GEN_1084 = _T_128 ? 4'h3 : _GEN_912; // @[FSM.scala 896:30 FSM.scala 900:21]
  wire [9:0] _GEN_1085 = gru_state == 4'h2 ? _GEN_1081 : _GEN_885; // @[FSM.scala 725:30]
  wire [6:0] _GEN_1086 = gru_state == 4'h2 ? _GEN_882 : _GEN_886; // @[FSM.scala 725:30]
  wire [2:0] _GEN_1087 = gru_state == 4'h2 ? _GEN_925 : _GEN_887; // @[FSM.scala 725:30]
  wire [9:0] _GEN_1088 = gru_state == 4'h2 ? _GEN_926 : _GEN_888; // @[FSM.scala 725:30]
  wire [5:0] _GEN_1089 = gru_state == 4'h2 ? _GEN_927 : _GEN_889; // @[FSM.scala 725:30]
  wire [11:0] _GEN_1090 = gru_state == 4'h2 ? _GEN_932 : _GEN_890; // @[FSM.scala 725:30]
  wire [7:0] _GEN_1091 = gru_state == 4'h2 ? _GEN_929 : _GEN_891; // @[FSM.scala 725:30]
  wire [1:0] _GEN_1092 = gru_state == 4'h2 ? _GEN_920 : _GEN_904; // @[FSM.scala 725:30]
  wire [3:0] _GEN_1093 = gru_state == 4'h2 ? _GEN_921 : _GEN_905; // @[FSM.scala 725:30]
  wire [5:0] _GEN_1094 = gru_state == 4'h2 ? _GEN_1079 : Rt_wrAddr; // @[FSM.scala 725:30 FSM.scala 86:36]
  wire [1:0] _GEN_1095 = gru_state == 4'h2 ? _GEN_923 : _GEN_907; // @[FSM.scala 725:30]
  wire [1:0] _GEN_1096 = gru_state == 4'h2 ? _GEN_924 : _GEN_908; // @[FSM.scala 725:30]
  wire [11:0] _GEN_1097 = gru_state == 4'h2 ? _GEN_930 : _GEN_909; // @[FSM.scala 725:30]
  wire [11:0] _GEN_1098 = gru_state == 4'h2 ? _GEN_931 : _GEN_910; // @[FSM.scala 725:30]
  wire [11:0] _GEN_1099 = gru_state == 4'h2 ? _GEN_999 : _GEN_892; // @[FSM.scala 725:30]
  wire [11:0] _GEN_1100 = gru_state == 4'h2 ? _GEN_1011 : _GEN_893; // @[FSM.scala 725:30]
  wire [11:0] _GEN_1101 = gru_state == 4'h2 ? _GEN_1022 : _GEN_894; // @[FSM.scala 725:30]
  wire [11:0] _GEN_1102 = gru_state == 4'h2 ? _GEN_1032 : _GEN_895; // @[FSM.scala 725:30]
  wire [11:0] _GEN_1103 = gru_state == 4'h2 ? _GEN_1041 : _GEN_896; // @[FSM.scala 725:30]
  wire [11:0] _GEN_1104 = gru_state == 4'h2 ? _GEN_1049 : _GEN_897; // @[FSM.scala 725:30]
  wire [11:0] _GEN_1105 = gru_state == 4'h2 ? _GEN_1056 : _GEN_898; // @[FSM.scala 725:30]
  wire [11:0] _GEN_1106 = gru_state == 4'h2 ? _GEN_1062 : _GEN_899; // @[FSM.scala 725:30]
  wire [11:0] _GEN_1107 = gru_state == 4'h2 ? _GEN_1067 : _GEN_900; // @[FSM.scala 725:30]
  wire [11:0] _GEN_1108 = gru_state == 4'h2 ? _GEN_1071 : _GEN_901; // @[FSM.scala 725:30]
  wire [11:0] _GEN_1109 = gru_state == 4'h2 ? _GEN_1074 : _GEN_902; // @[FSM.scala 725:30]
  wire [11:0] _GEN_1110 = gru_state == 4'h2 ? _GEN_1076 : _GEN_903; // @[FSM.scala 725:30]
  wire  _GEN_1111 = gru_state == 4'h2 ? _GEN_1083 : Rt_wrEna; // @[FSM.scala 725:30 FSM.scala 85:36]
  wire [3:0] _GEN_1112 = gru_state == 4'h2 ? _GEN_1084 : _GEN_912; // @[FSM.scala 725:30]
  wire [9:0] _GEN_1113 = count != 10'h20e ? _count_T_1 : _GEN_1085; // @[FSM.scala 906:30 FSM.scala 907:17]
  wire [2:0] _GEN_1115 = _T_3 ? 3'h4 : _GEN_1087; // @[FSM.scala 916:28 FSM.scala 918:35]
  wire [9:0] _GEN_1116 = _T_3 ? 10'h1ff : _GEN_1088; // @[FSM.scala 916:28 FSM.scala 919:33]
  wire [5:0] _GEN_1117 = _T_3 ? 6'h15 : _GEN_1089; // @[FSM.scala 916:28 FSM.scala 920:35]
  wire [11:0] _GEN_1118 = _T_3 ? 12'h800 : _GEN_1090; // @[FSM.scala 916:28 FSM.scala 921:32]
  wire [7:0] _GEN_1119 = _T_3 ? 8'h40 : _GEN_1091; // @[FSM.scala 916:28 FSM.scala 922:41]
  wire [1:0] _GEN_1120 = _T_3 ? 2'h0 : _GEN_1092; // @[FSM.scala 916:28 FSM.scala 925:30]
  wire [3:0] _GEN_1121 = _T_3 ? 4'h0 : _GEN_1093; // @[FSM.scala 916:28 FSM.scala 926:26]
  wire [5:0] _GEN_1122 = _T_3 ? 6'h0 : WhXt_wrAddr; // @[FSM.scala 916:28 FSM.scala 929:23 FSM.scala 89:36]
  wire [1:0] _GEN_1123 = _T_3 ? 2'h0 : _GEN_1095; // @[FSM.scala 916:28 FSM.scala 930:24]
  wire [1:0] _GEN_1124 = _T_3 ? 2'h0 : _GEN_1096; // @[FSM.scala 916:28 FSM.scala 931:27]
  wire [2:0] _GEN_1125 = _T_39 ? 3'h4 : _GEN_1115; // @[FSM.scala 935:48 FSM.scala 936:35]
  wire [9:0] _GEN_1126 = _T_39 ? 10'h1ff : _GEN_1116; // @[FSM.scala 935:48 FSM.scala 937:33]
  wire [5:0] _GEN_1127 = _T_39 ? 6'h15 : _GEN_1117; // @[FSM.scala 935:48 FSM.scala 938:35]
  wire [11:0] _GEN_1128 = _T_39 ? {{1'd0}, PEArray_ctrl_2_mask[11:1]} : _GEN_1118; // @[FSM.scala 935:48 FSM.scala 939:32]
  wire [7:0] _GEN_1129 = _T_39 ? 8'h40 : _GEN_1119; // @[FSM.scala 935:48 FSM.scala 940:41]
  wire [11:0] _GEN_1130 = _T_40 ? 12'h0 : _GEN_1097; // @[FSM.scala 942:29 FSM.scala 944:34]
  wire [11:0] _GEN_1131 = _T_40 ? 12'h0 : _GEN_1098; // @[FSM.scala 942:29 FSM.scala 944:34]
  wire [11:0] _GEN_1132 = _T_40 ? 12'h0 : _GEN_1128; // @[FSM.scala 942:29 FSM.scala 944:34]
  wire [11:0] _GEN_1133 = _T_5 ? _L1_rd_addr_0_T_1 : _GEN_1099; // @[FSM.scala 949:28 FSM.scala 951:27]
  wire [11:0] _GEN_1134 = _T_48 ? _L1_rd_addr_0_T_1 : _GEN_1133; // @[FSM.scala 954:28 FSM.scala 956:27]
  wire [11:0] _GEN_1135 = _T_48 ? _L1_rd_addr_1_T_1 : _GEN_1100; // @[FSM.scala 954:28 FSM.scala 956:27]
  wire [11:0] _GEN_1136 = _T_49 ? _L1_rd_addr_0_T_1 : _GEN_1134; // @[FSM.scala 959:28 FSM.scala 961:27]
  wire [11:0] _GEN_1137 = _T_49 ? _L1_rd_addr_1_T_1 : _GEN_1135; // @[FSM.scala 959:28 FSM.scala 961:27]
  wire [11:0] _GEN_1138 = _T_49 ? _L1_rd_addr_2_T_1 : _GEN_1101; // @[FSM.scala 959:28 FSM.scala 961:27]
  wire [11:0] _GEN_1139 = _T_21 ? _L1_rd_addr_0_T_1 : _GEN_1136; // @[FSM.scala 964:28 FSM.scala 966:27]
  wire [11:0] _GEN_1140 = _T_21 ? _L1_rd_addr_1_T_1 : _GEN_1137; // @[FSM.scala 964:28 FSM.scala 966:27]
  wire [11:0] _GEN_1141 = _T_21 ? _L1_rd_addr_2_T_1 : _GEN_1138; // @[FSM.scala 964:28 FSM.scala 966:27]
  wire [11:0] _GEN_1142 = _T_21 ? _L1_rd_addr_3_T_1 : _GEN_1102; // @[FSM.scala 964:28 FSM.scala 966:27]
  wire [11:0] _GEN_1143 = _T_51 ? _L1_rd_addr_0_T_1 : _GEN_1139; // @[FSM.scala 969:28 FSM.scala 971:27]
  wire [11:0] _GEN_1144 = _T_51 ? _L1_rd_addr_1_T_1 : _GEN_1140; // @[FSM.scala 969:28 FSM.scala 971:27]
  wire [11:0] _GEN_1145 = _T_51 ? _L1_rd_addr_2_T_1 : _GEN_1141; // @[FSM.scala 969:28 FSM.scala 971:27]
  wire [11:0] _GEN_1146 = _T_51 ? _L1_rd_addr_3_T_1 : _GEN_1142; // @[FSM.scala 969:28 FSM.scala 971:27]
  wire [11:0] _GEN_1147 = _T_51 ? _L1_rd_addr_4_T_1 : _GEN_1103; // @[FSM.scala 969:28 FSM.scala 971:27]
  wire [11:0] _GEN_1148 = _T_52 ? _L1_rd_addr_0_T_1 : _GEN_1143; // @[FSM.scala 974:28 FSM.scala 976:27]
  wire [11:0] _GEN_1149 = _T_52 ? _L1_rd_addr_1_T_1 : _GEN_1144; // @[FSM.scala 974:28 FSM.scala 976:27]
  wire [11:0] _GEN_1150 = _T_52 ? _L1_rd_addr_2_T_1 : _GEN_1145; // @[FSM.scala 974:28 FSM.scala 976:27]
  wire [11:0] _GEN_1151 = _T_52 ? _L1_rd_addr_3_T_1 : _GEN_1146; // @[FSM.scala 974:28 FSM.scala 976:27]
  wire [11:0] _GEN_1152 = _T_52 ? _L1_rd_addr_4_T_1 : _GEN_1147; // @[FSM.scala 974:28 FSM.scala 976:27]
  wire [11:0] _GEN_1153 = _T_52 ? _L1_rd_addr_5_T_1 : _GEN_1104; // @[FSM.scala 974:28 FSM.scala 976:27]
  wire [11:0] _GEN_1154 = _T_53 ? _L1_rd_addr_0_T_1 : _GEN_1148; // @[FSM.scala 979:28 FSM.scala 981:27]
  wire [11:0] _GEN_1155 = _T_53 ? _L1_rd_addr_1_T_1 : _GEN_1149; // @[FSM.scala 979:28 FSM.scala 981:27]
  wire [11:0] _GEN_1156 = _T_53 ? _L1_rd_addr_2_T_1 : _GEN_1150; // @[FSM.scala 979:28 FSM.scala 981:27]
  wire [11:0] _GEN_1157 = _T_53 ? _L1_rd_addr_3_T_1 : _GEN_1151; // @[FSM.scala 979:28 FSM.scala 981:27]
  wire [11:0] _GEN_1158 = _T_53 ? _L1_rd_addr_4_T_1 : _GEN_1152; // @[FSM.scala 979:28 FSM.scala 981:27]
  wire [11:0] _GEN_1159 = _T_53 ? _L1_rd_addr_5_T_1 : _GEN_1153; // @[FSM.scala 979:28 FSM.scala 981:27]
  wire [11:0] _GEN_1160 = _T_53 ? _L1_rd_addr_6_T_1 : _GEN_1105; // @[FSM.scala 979:28 FSM.scala 981:27]
  wire [11:0] _GEN_1161 = _T_54 ? _L1_rd_addr_0_T_1 : _GEN_1154; // @[FSM.scala 984:28 FSM.scala 986:27]
  wire [11:0] _GEN_1162 = _T_54 ? _L1_rd_addr_1_T_1 : _GEN_1155; // @[FSM.scala 984:28 FSM.scala 986:27]
  wire [11:0] _GEN_1163 = _T_54 ? _L1_rd_addr_2_T_1 : _GEN_1156; // @[FSM.scala 984:28 FSM.scala 986:27]
  wire [11:0] _GEN_1164 = _T_54 ? _L1_rd_addr_3_T_1 : _GEN_1157; // @[FSM.scala 984:28 FSM.scala 986:27]
  wire [11:0] _GEN_1165 = _T_54 ? _L1_rd_addr_4_T_1 : _GEN_1158; // @[FSM.scala 984:28 FSM.scala 986:27]
  wire [11:0] _GEN_1166 = _T_54 ? _L1_rd_addr_5_T_1 : _GEN_1159; // @[FSM.scala 984:28 FSM.scala 986:27]
  wire [11:0] _GEN_1167 = _T_54 ? _L1_rd_addr_6_T_1 : _GEN_1160; // @[FSM.scala 984:28 FSM.scala 986:27]
  wire [11:0] _GEN_1168 = _T_54 ? _L1_rd_addr_7_T_1 : _GEN_1106; // @[FSM.scala 984:28 FSM.scala 986:27]
  wire [11:0] _GEN_1169 = _T_55 ? _L1_rd_addr_0_T_1 : _GEN_1161; // @[FSM.scala 989:28 FSM.scala 991:27]
  wire [11:0] _GEN_1170 = _T_55 ? _L1_rd_addr_1_T_1 : _GEN_1162; // @[FSM.scala 989:28 FSM.scala 991:27]
  wire [11:0] _GEN_1171 = _T_55 ? _L1_rd_addr_2_T_1 : _GEN_1163; // @[FSM.scala 989:28 FSM.scala 991:27]
  wire [11:0] _GEN_1172 = _T_55 ? _L1_rd_addr_3_T_1 : _GEN_1164; // @[FSM.scala 989:28 FSM.scala 991:27]
  wire [11:0] _GEN_1173 = _T_55 ? _L1_rd_addr_4_T_1 : _GEN_1165; // @[FSM.scala 989:28 FSM.scala 991:27]
  wire [11:0] _GEN_1174 = _T_55 ? _L1_rd_addr_5_T_1 : _GEN_1166; // @[FSM.scala 989:28 FSM.scala 991:27]
  wire [11:0] _GEN_1175 = _T_55 ? _L1_rd_addr_6_T_1 : _GEN_1167; // @[FSM.scala 989:28 FSM.scala 991:27]
  wire [11:0] _GEN_1176 = _T_55 ? _L1_rd_addr_7_T_1 : _GEN_1168; // @[FSM.scala 989:28 FSM.scala 991:27]
  wire [11:0] _GEN_1177 = _T_55 ? _L1_rd_addr_8_T_1 : _GEN_1107; // @[FSM.scala 989:28 FSM.scala 991:27]
  wire [11:0] _GEN_1178 = _T_56 ? _L1_rd_addr_0_T_1 : _GEN_1169; // @[FSM.scala 994:29 FSM.scala 996:27]
  wire [11:0] _GEN_1179 = _T_56 ? _L1_rd_addr_1_T_1 : _GEN_1170; // @[FSM.scala 994:29 FSM.scala 996:27]
  wire [11:0] _GEN_1180 = _T_56 ? _L1_rd_addr_2_T_1 : _GEN_1171; // @[FSM.scala 994:29 FSM.scala 996:27]
  wire [11:0] _GEN_1181 = _T_56 ? _L1_rd_addr_3_T_1 : _GEN_1172; // @[FSM.scala 994:29 FSM.scala 996:27]
  wire [11:0] _GEN_1182 = _T_56 ? _L1_rd_addr_4_T_1 : _GEN_1173; // @[FSM.scala 994:29 FSM.scala 996:27]
  wire [11:0] _GEN_1183 = _T_56 ? _L1_rd_addr_5_T_1 : _GEN_1174; // @[FSM.scala 994:29 FSM.scala 996:27]
  wire [11:0] _GEN_1184 = _T_56 ? _L1_rd_addr_6_T_1 : _GEN_1175; // @[FSM.scala 994:29 FSM.scala 996:27]
  wire [11:0] _GEN_1185 = _T_56 ? _L1_rd_addr_7_T_1 : _GEN_1176; // @[FSM.scala 994:29 FSM.scala 996:27]
  wire [11:0] _GEN_1186 = _T_56 ? _L1_rd_addr_8_T_1 : _GEN_1177; // @[FSM.scala 994:29 FSM.scala 996:27]
  wire [11:0] _GEN_1187 = _T_56 ? _L1_rd_addr_9_T_1 : _GEN_1108; // @[FSM.scala 994:29 FSM.scala 996:27]
  wire [11:0] _GEN_1188 = _T_57 ? _L1_rd_addr_0_T_1 : _GEN_1178; // @[FSM.scala 999:29 FSM.scala 1001:27]
  wire [11:0] _GEN_1189 = _T_57 ? _L1_rd_addr_1_T_1 : _GEN_1179; // @[FSM.scala 999:29 FSM.scala 1001:27]
  wire [11:0] _GEN_1190 = _T_57 ? _L1_rd_addr_2_T_1 : _GEN_1180; // @[FSM.scala 999:29 FSM.scala 1001:27]
  wire [11:0] _GEN_1191 = _T_57 ? _L1_rd_addr_3_T_1 : _GEN_1181; // @[FSM.scala 999:29 FSM.scala 1001:27]
  wire [11:0] _GEN_1192 = _T_57 ? _L1_rd_addr_4_T_1 : _GEN_1182; // @[FSM.scala 999:29 FSM.scala 1001:27]
  wire [11:0] _GEN_1193 = _T_57 ? _L1_rd_addr_5_T_1 : _GEN_1183; // @[FSM.scala 999:29 FSM.scala 1001:27]
  wire [11:0] _GEN_1194 = _T_57 ? _L1_rd_addr_6_T_1 : _GEN_1184; // @[FSM.scala 999:29 FSM.scala 1001:27]
  wire [11:0] _GEN_1195 = _T_57 ? _L1_rd_addr_7_T_1 : _GEN_1185; // @[FSM.scala 999:29 FSM.scala 1001:27]
  wire [11:0] _GEN_1196 = _T_57 ? _L1_rd_addr_8_T_1 : _GEN_1186; // @[FSM.scala 999:29 FSM.scala 1001:27]
  wire [11:0] _GEN_1197 = _T_57 ? _L1_rd_addr_9_T_1 : _GEN_1187; // @[FSM.scala 999:29 FSM.scala 1001:27]
  wire [11:0] _GEN_1198 = _T_57 ? _L1_rd_addr_10_T_1 : _GEN_1109; // @[FSM.scala 999:29 FSM.scala 1001:27]
  wire [11:0] _GEN_1199 = _T_110 & count <= 10'h1ff ? _L1_rd_addr_0_T_1 : _GEN_1188; // @[FSM.scala 1004:50 FSM.scala 1006:27]
  wire [11:0] _GEN_1200 = _T_110 & count <= 10'h1ff ? _L1_rd_addr_1_T_1 : _GEN_1189; // @[FSM.scala 1004:50 FSM.scala 1006:27]
  wire [11:0] _GEN_1201 = _T_110 & count <= 10'h1ff ? _L1_rd_addr_2_T_1 : _GEN_1190; // @[FSM.scala 1004:50 FSM.scala 1006:27]
  wire [11:0] _GEN_1202 = _T_110 & count <= 10'h1ff ? _L1_rd_addr_3_T_1 : _GEN_1191; // @[FSM.scala 1004:50 FSM.scala 1006:27]
  wire [11:0] _GEN_1203 = _T_110 & count <= 10'h1ff ? _L1_rd_addr_4_T_1 : _GEN_1192; // @[FSM.scala 1004:50 FSM.scala 1006:27]
  wire [11:0] _GEN_1204 = _T_110 & count <= 10'h1ff ? _L1_rd_addr_5_T_1 : _GEN_1193; // @[FSM.scala 1004:50 FSM.scala 1006:27]
  wire [11:0] _GEN_1205 = _T_110 & count <= 10'h1ff ? _L1_rd_addr_6_T_1 : _GEN_1194; // @[FSM.scala 1004:50 FSM.scala 1006:27]
  wire [11:0] _GEN_1206 = _T_110 & count <= 10'h1ff ? _L1_rd_addr_7_T_1 : _GEN_1195; // @[FSM.scala 1004:50 FSM.scala 1006:27]
  wire [11:0] _GEN_1207 = _T_110 & count <= 10'h1ff ? _L1_rd_addr_8_T_1 : _GEN_1196; // @[FSM.scala 1004:50 FSM.scala 1006:27]
  wire [11:0] _GEN_1208 = _T_110 & count <= 10'h1ff ? _L1_rd_addr_9_T_1 : _GEN_1197; // @[FSM.scala 1004:50 FSM.scala 1006:27]
  wire [11:0] _GEN_1209 = _T_110 & count <= 10'h1ff ? _L1_rd_addr_10_T_1 : _GEN_1198; // @[FSM.scala 1004:50 FSM.scala 1006:27]
  wire [11:0] _GEN_1210 = _T_110 & count <= 10'h1ff ? _L1_rd_addr_11_T_1 : _GEN_1110; // @[FSM.scala 1004:50 FSM.scala 1006:27]
  wire [11:0] _GEN_1211 = count == 10'h200 ? _L1_rd_addr_1_T_1 : _GEN_1200; // @[FSM.scala 1009:30 FSM.scala 1011:27]
  wire [11:0] _GEN_1212 = count == 10'h200 ? _L1_rd_addr_2_T_1 : _GEN_1201; // @[FSM.scala 1009:30 FSM.scala 1011:27]
  wire [11:0] _GEN_1213 = count == 10'h200 ? _L1_rd_addr_3_T_1 : _GEN_1202; // @[FSM.scala 1009:30 FSM.scala 1011:27]
  wire [11:0] _GEN_1214 = count == 10'h200 ? _L1_rd_addr_4_T_1 : _GEN_1203; // @[FSM.scala 1009:30 FSM.scala 1011:27]
  wire [11:0] _GEN_1215 = count == 10'h200 ? _L1_rd_addr_5_T_1 : _GEN_1204; // @[FSM.scala 1009:30 FSM.scala 1011:27]
  wire [11:0] _GEN_1216 = count == 10'h200 ? _L1_rd_addr_6_T_1 : _GEN_1205; // @[FSM.scala 1009:30 FSM.scala 1011:27]
  wire [11:0] _GEN_1217 = count == 10'h200 ? _L1_rd_addr_7_T_1 : _GEN_1206; // @[FSM.scala 1009:30 FSM.scala 1011:27]
  wire [11:0] _GEN_1218 = count == 10'h200 ? _L1_rd_addr_8_T_1 : _GEN_1207; // @[FSM.scala 1009:30 FSM.scala 1011:27]
  wire [11:0] _GEN_1219 = count == 10'h200 ? _L1_rd_addr_9_T_1 : _GEN_1208; // @[FSM.scala 1009:30 FSM.scala 1011:27]
  wire [11:0] _GEN_1220 = count == 10'h200 ? _L1_rd_addr_10_T_1 : _GEN_1209; // @[FSM.scala 1009:30 FSM.scala 1011:27]
  wire [11:0] _GEN_1221 = count == 10'h200 ? _L1_rd_addr_11_T_1 : _GEN_1210; // @[FSM.scala 1009:30 FSM.scala 1011:27]
  wire [11:0] _GEN_1222 = count == 10'h201 ? _L1_rd_addr_2_T_1 : _GEN_1212; // @[FSM.scala 1014:30 FSM.scala 1016:27]
  wire [11:0] _GEN_1223 = count == 10'h201 ? _L1_rd_addr_3_T_1 : _GEN_1213; // @[FSM.scala 1014:30 FSM.scala 1016:27]
  wire [11:0] _GEN_1224 = count == 10'h201 ? _L1_rd_addr_4_T_1 : _GEN_1214; // @[FSM.scala 1014:30 FSM.scala 1016:27]
  wire [11:0] _GEN_1225 = count == 10'h201 ? _L1_rd_addr_5_T_1 : _GEN_1215; // @[FSM.scala 1014:30 FSM.scala 1016:27]
  wire [11:0] _GEN_1226 = count == 10'h201 ? _L1_rd_addr_6_T_1 : _GEN_1216; // @[FSM.scala 1014:30 FSM.scala 1016:27]
  wire [11:0] _GEN_1227 = count == 10'h201 ? _L1_rd_addr_7_T_1 : _GEN_1217; // @[FSM.scala 1014:30 FSM.scala 1016:27]
  wire [11:0] _GEN_1228 = count == 10'h201 ? _L1_rd_addr_8_T_1 : _GEN_1218; // @[FSM.scala 1014:30 FSM.scala 1016:27]
  wire [11:0] _GEN_1229 = count == 10'h201 ? _L1_rd_addr_9_T_1 : _GEN_1219; // @[FSM.scala 1014:30 FSM.scala 1016:27]
  wire [11:0] _GEN_1230 = count == 10'h201 ? _L1_rd_addr_10_T_1 : _GEN_1220; // @[FSM.scala 1014:30 FSM.scala 1016:27]
  wire [11:0] _GEN_1231 = count == 10'h201 ? _L1_rd_addr_11_T_1 : _GEN_1221; // @[FSM.scala 1014:30 FSM.scala 1016:27]
  wire [11:0] _GEN_1232 = count == 10'h202 ? _L1_rd_addr_3_T_1 : _GEN_1223; // @[FSM.scala 1019:30 FSM.scala 1021:27]
  wire [11:0] _GEN_1233 = count == 10'h202 ? _L1_rd_addr_4_T_1 : _GEN_1224; // @[FSM.scala 1019:30 FSM.scala 1021:27]
  wire [11:0] _GEN_1234 = count == 10'h202 ? _L1_rd_addr_5_T_1 : _GEN_1225; // @[FSM.scala 1019:30 FSM.scala 1021:27]
  wire [11:0] _GEN_1235 = count == 10'h202 ? _L1_rd_addr_6_T_1 : _GEN_1226; // @[FSM.scala 1019:30 FSM.scala 1021:27]
  wire [11:0] _GEN_1236 = count == 10'h202 ? _L1_rd_addr_7_T_1 : _GEN_1227; // @[FSM.scala 1019:30 FSM.scala 1021:27]
  wire [11:0] _GEN_1237 = count == 10'h202 ? _L1_rd_addr_8_T_1 : _GEN_1228; // @[FSM.scala 1019:30 FSM.scala 1021:27]
  wire [11:0] _GEN_1238 = count == 10'h202 ? _L1_rd_addr_9_T_1 : _GEN_1229; // @[FSM.scala 1019:30 FSM.scala 1021:27]
  wire [11:0] _GEN_1239 = count == 10'h202 ? _L1_rd_addr_10_T_1 : _GEN_1230; // @[FSM.scala 1019:30 FSM.scala 1021:27]
  wire [11:0] _GEN_1240 = count == 10'h202 ? _L1_rd_addr_11_T_1 : _GEN_1231; // @[FSM.scala 1019:30 FSM.scala 1021:27]
  wire [11:0] _GEN_1241 = count == 10'h203 ? _L1_rd_addr_4_T_1 : _GEN_1233; // @[FSM.scala 1024:30 FSM.scala 1026:27]
  wire [11:0] _GEN_1242 = count == 10'h203 ? _L1_rd_addr_5_T_1 : _GEN_1234; // @[FSM.scala 1024:30 FSM.scala 1026:27]
  wire [11:0] _GEN_1243 = count == 10'h203 ? _L1_rd_addr_6_T_1 : _GEN_1235; // @[FSM.scala 1024:30 FSM.scala 1026:27]
  wire [11:0] _GEN_1244 = count == 10'h203 ? _L1_rd_addr_7_T_1 : _GEN_1236; // @[FSM.scala 1024:30 FSM.scala 1026:27]
  wire [11:0] _GEN_1245 = count == 10'h203 ? _L1_rd_addr_8_T_1 : _GEN_1237; // @[FSM.scala 1024:30 FSM.scala 1026:27]
  wire [11:0] _GEN_1246 = count == 10'h203 ? _L1_rd_addr_9_T_1 : _GEN_1238; // @[FSM.scala 1024:30 FSM.scala 1026:27]
  wire [11:0] _GEN_1247 = count == 10'h203 ? _L1_rd_addr_10_T_1 : _GEN_1239; // @[FSM.scala 1024:30 FSM.scala 1026:27]
  wire [11:0] _GEN_1248 = count == 10'h203 ? _L1_rd_addr_11_T_1 : _GEN_1240; // @[FSM.scala 1024:30 FSM.scala 1026:27]
  wire [11:0] _GEN_1249 = count == 10'h204 ? _L1_rd_addr_5_T_1 : _GEN_1242; // @[FSM.scala 1029:30 FSM.scala 1031:27]
  wire [11:0] _GEN_1250 = count == 10'h204 ? _L1_rd_addr_6_T_1 : _GEN_1243; // @[FSM.scala 1029:30 FSM.scala 1031:27]
  wire [11:0] _GEN_1251 = count == 10'h204 ? _L1_rd_addr_7_T_1 : _GEN_1244; // @[FSM.scala 1029:30 FSM.scala 1031:27]
  wire [11:0] _GEN_1252 = count == 10'h204 ? _L1_rd_addr_8_T_1 : _GEN_1245; // @[FSM.scala 1029:30 FSM.scala 1031:27]
  wire [11:0] _GEN_1253 = count == 10'h204 ? _L1_rd_addr_9_T_1 : _GEN_1246; // @[FSM.scala 1029:30 FSM.scala 1031:27]
  wire [11:0] _GEN_1254 = count == 10'h204 ? _L1_rd_addr_10_T_1 : _GEN_1247; // @[FSM.scala 1029:30 FSM.scala 1031:27]
  wire [11:0] _GEN_1255 = count == 10'h204 ? _L1_rd_addr_11_T_1 : _GEN_1248; // @[FSM.scala 1029:30 FSM.scala 1031:27]
  wire [11:0] _GEN_1256 = count == 10'h205 ? _L1_rd_addr_6_T_1 : _GEN_1250; // @[FSM.scala 1034:30 FSM.scala 1036:27]
  wire [11:0] _GEN_1257 = count == 10'h205 ? _L1_rd_addr_7_T_1 : _GEN_1251; // @[FSM.scala 1034:30 FSM.scala 1036:27]
  wire [11:0] _GEN_1258 = count == 10'h205 ? _L1_rd_addr_8_T_1 : _GEN_1252; // @[FSM.scala 1034:30 FSM.scala 1036:27]
  wire [11:0] _GEN_1259 = count == 10'h205 ? _L1_rd_addr_9_T_1 : _GEN_1253; // @[FSM.scala 1034:30 FSM.scala 1036:27]
  wire [11:0] _GEN_1260 = count == 10'h205 ? _L1_rd_addr_10_T_1 : _GEN_1254; // @[FSM.scala 1034:30 FSM.scala 1036:27]
  wire [11:0] _GEN_1261 = count == 10'h205 ? _L1_rd_addr_11_T_1 : _GEN_1255; // @[FSM.scala 1034:30 FSM.scala 1036:27]
  wire [11:0] _GEN_1262 = count == 10'h206 ? _L1_rd_addr_7_T_1 : _GEN_1257; // @[FSM.scala 1039:30 FSM.scala 1041:27]
  wire [11:0] _GEN_1263 = count == 10'h206 ? _L1_rd_addr_8_T_1 : _GEN_1258; // @[FSM.scala 1039:30 FSM.scala 1041:27]
  wire [11:0] _GEN_1264 = count == 10'h206 ? _L1_rd_addr_9_T_1 : _GEN_1259; // @[FSM.scala 1039:30 FSM.scala 1041:27]
  wire [11:0] _GEN_1265 = count == 10'h206 ? _L1_rd_addr_10_T_1 : _GEN_1260; // @[FSM.scala 1039:30 FSM.scala 1041:27]
  wire [11:0] _GEN_1266 = count == 10'h206 ? _L1_rd_addr_11_T_1 : _GEN_1261; // @[FSM.scala 1039:30 FSM.scala 1041:27]
  wire [11:0] _GEN_1267 = count == 10'h207 ? _L1_rd_addr_8_T_1 : _GEN_1263; // @[FSM.scala 1044:30 FSM.scala 1046:27]
  wire [11:0] _GEN_1268 = count == 10'h207 ? _L1_rd_addr_9_T_1 : _GEN_1264; // @[FSM.scala 1044:30 FSM.scala 1046:27]
  wire [11:0] _GEN_1269 = count == 10'h207 ? _L1_rd_addr_10_T_1 : _GEN_1265; // @[FSM.scala 1044:30 FSM.scala 1046:27]
  wire [11:0] _GEN_1270 = count == 10'h207 ? _L1_rd_addr_11_T_1 : _GEN_1266; // @[FSM.scala 1044:30 FSM.scala 1046:27]
  wire [11:0] _GEN_1271 = count == 10'h208 ? _L1_rd_addr_9_T_1 : _GEN_1268; // @[FSM.scala 1049:30 FSM.scala 1051:27]
  wire [11:0] _GEN_1272 = count == 10'h208 ? _L1_rd_addr_10_T_1 : _GEN_1269; // @[FSM.scala 1049:30 FSM.scala 1051:27]
  wire [11:0] _GEN_1273 = count == 10'h208 ? _L1_rd_addr_11_T_1 : _GEN_1270; // @[FSM.scala 1049:30 FSM.scala 1051:27]
  wire [11:0] _GEN_1274 = count == 10'h209 ? _L1_rd_addr_10_T_1 : _GEN_1272; // @[FSM.scala 1054:30 FSM.scala 1056:27]
  wire [11:0] _GEN_1275 = count == 10'h209 ? _L1_rd_addr_11_T_1 : _GEN_1273; // @[FSM.scala 1054:30 FSM.scala 1056:27]
  wire [11:0] _GEN_1276 = count == 10'h20a ? _L1_rd_addr_11_T_1 : _GEN_1275; // @[FSM.scala 1059:30 FSM.scala 1061:27]
  wire [5:0] _WhXt_wrAddr_T_1 = WhXt_wrAddr + 6'h1; // @[FSM.scala 1071:42]
  wire [5:0] _GEN_1277 = _T_127 ? 6'h0 : _WhXt_wrAddr_T_1; // @[FSM.scala 1066:33 FSM.scala 1067:25 FSM.scala 1071:27]
  wire [5:0] _GEN_1279 = _T_124 & count <= 10'h20d ? _GEN_1277 : _GEN_1122; // @[FSM.scala 1065:50]
  wire  _GEN_1280 = _T_124 & count <= 10'h20d | WhXt_wrEna; // @[FSM.scala 1065:50 FSM.scala 88:36]
  wire [9:0] _GEN_1281 = count == 10'h20e ? 10'h0 : _GEN_1113; // @[FSM.scala 1076:30 FSM.scala 1077:17]
  wire [6:0] _GEN_1282 = count == 10'h20e ? 7'h0 : _GEN_702; // @[FSM.scala 1076:30 FSM.scala 1078:18]
  wire  _GEN_1283 = count == 10'h20e ? 1'h0 : _GEN_1280; // @[FSM.scala 1076:30 FSM.scala 1079:22]
  wire [3:0] _GEN_1284 = count == 10'h20e ? 4'h4 : _GEN_1112; // @[FSM.scala 1076:30 FSM.scala 1080:21]
  wire [9:0] _GEN_1285 = gru_state == 4'h3 ? _GEN_1281 : _GEN_1085; // @[FSM.scala 905:30]
  wire [6:0] _GEN_1286 = gru_state == 4'h3 ? _GEN_1282 : _GEN_1086; // @[FSM.scala 905:30]
  wire [2:0] _GEN_1287 = gru_state == 4'h3 ? _GEN_1125 : _GEN_1087; // @[FSM.scala 905:30]
  wire [9:0] _GEN_1288 = gru_state == 4'h3 ? _GEN_1126 : _GEN_1088; // @[FSM.scala 905:30]
  wire [5:0] _GEN_1289 = gru_state == 4'h3 ? _GEN_1127 : _GEN_1089; // @[FSM.scala 905:30]
  wire [11:0] _GEN_1290 = gru_state == 4'h3 ? _GEN_1132 : _GEN_1090; // @[FSM.scala 905:30]
  wire [7:0] _GEN_1291 = gru_state == 4'h3 ? _GEN_1129 : _GEN_1091; // @[FSM.scala 905:30]
  wire [1:0] _GEN_1292 = gru_state == 4'h3 ? _GEN_1120 : _GEN_1092; // @[FSM.scala 905:30]
  wire [3:0] _GEN_1293 = gru_state == 4'h3 ? _GEN_1121 : _GEN_1093; // @[FSM.scala 905:30]
  wire [5:0] _GEN_1294 = gru_state == 4'h3 ? _GEN_1279 : WhXt_wrAddr; // @[FSM.scala 905:30 FSM.scala 89:36]
  wire [1:0] _GEN_1295 = gru_state == 4'h3 ? _GEN_1123 : _GEN_1095; // @[FSM.scala 905:30]
  wire [1:0] _GEN_1296 = gru_state == 4'h3 ? _GEN_1124 : _GEN_1096; // @[FSM.scala 905:30]
  wire [11:0] _GEN_1297 = gru_state == 4'h3 ? _GEN_1130 : _GEN_1097; // @[FSM.scala 905:30]
  wire [11:0] _GEN_1298 = gru_state == 4'h3 ? _GEN_1131 : _GEN_1098; // @[FSM.scala 905:30]
  wire [11:0] _GEN_1299 = gru_state == 4'h3 ? _GEN_1199 : _GEN_1099; // @[FSM.scala 905:30]
  wire [11:0] _GEN_1300 = gru_state == 4'h3 ? _GEN_1211 : _GEN_1100; // @[FSM.scala 905:30]
  wire [11:0] _GEN_1301 = gru_state == 4'h3 ? _GEN_1222 : _GEN_1101; // @[FSM.scala 905:30]
  wire [11:0] _GEN_1302 = gru_state == 4'h3 ? _GEN_1232 : _GEN_1102; // @[FSM.scala 905:30]
  wire [11:0] _GEN_1303 = gru_state == 4'h3 ? _GEN_1241 : _GEN_1103; // @[FSM.scala 905:30]
  wire [11:0] _GEN_1304 = gru_state == 4'h3 ? _GEN_1249 : _GEN_1104; // @[FSM.scala 905:30]
  wire [11:0] _GEN_1305 = gru_state == 4'h3 ? _GEN_1256 : _GEN_1105; // @[FSM.scala 905:30]
  wire [11:0] _GEN_1306 = gru_state == 4'h3 ? _GEN_1262 : _GEN_1106; // @[FSM.scala 905:30]
  wire [11:0] _GEN_1307 = gru_state == 4'h3 ? _GEN_1267 : _GEN_1107; // @[FSM.scala 905:30]
  wire [11:0] _GEN_1308 = gru_state == 4'h3 ? _GEN_1271 : _GEN_1108; // @[FSM.scala 905:30]
  wire [11:0] _GEN_1309 = gru_state == 4'h3 ? _GEN_1274 : _GEN_1109; // @[FSM.scala 905:30]
  wire [11:0] _GEN_1310 = gru_state == 4'h3 ? _GEN_1276 : _GEN_1110; // @[FSM.scala 905:30]
  wire  _GEN_1311 = gru_state == 4'h3 ? _GEN_1283 : WhXt_wrEna; // @[FSM.scala 905:30 FSM.scala 88:36]
  wire [3:0] _GEN_1312 = gru_state == 4'h3 ? _GEN_1284 : _GEN_1112; // @[FSM.scala 905:30]
  wire  _T_206 = count != 10'h18e; // @[FSM.scala 1086:20]
  wire [9:0] _GEN_1313 = count != 10'h18e ? _count_T_1 : _GEN_1285; // @[FSM.scala 1086:30 FSM.scala 1087:17]
  wire [2:0] _GEN_1315 = _T_3 ? 3'h4 : _GEN_1287; // @[FSM.scala 1097:28 FSM.scala 1099:35]
  wire [9:0] _GEN_1316 = _T_3 ? 10'h17f : _GEN_1288; // @[FSM.scala 1097:28 FSM.scala 1100:33]
  wire [5:0] _GEN_1317 = _T_3 ? 6'hf : _GEN_1289; // @[FSM.scala 1097:28 FSM.scala 1101:35]
  wire [11:0] _GEN_1318 = _T_3 ? 12'h800 : _GEN_1290; // @[FSM.scala 1097:28 FSM.scala 1102:32]
  wire [7:0] _GEN_1319 = _T_3 ? 8'h40 : _GEN_1291; // @[FSM.scala 1097:28 FSM.scala 1103:41]
  wire [1:0] _GEN_1320 = _T_3 ? 2'h0 : _GEN_1292; // @[FSM.scala 1097:28 FSM.scala 1106:30]
  wire [3:0] _GEN_1321 = _T_3 ? 4'h0 : _GEN_1293; // @[FSM.scala 1097:28 FSM.scala 1107:26]
  wire [5:0] _GEN_1322 = _T_3 ? 6'h0 : Uhht_1_wrAddr; // @[FSM.scala 1097:28 FSM.scala 1110:25 FSM.scala 92:36]
  wire [1:0] _GEN_1323 = _T_3 ? 2'h0 : _GEN_1295; // @[FSM.scala 1097:28 FSM.scala 1111:24]
  wire [1:0] _GEN_1324 = _T_3 ? 2'h0 : _GEN_1296; // @[FSM.scala 1097:28 FSM.scala 1112:27]
  wire [2:0] _GEN_1325 = _T_39 ? 3'h4 : _GEN_1315; // @[FSM.scala 1116:48 FSM.scala 1117:35]
  wire [9:0] _GEN_1326 = _T_39 ? 10'h17f : _GEN_1316; // @[FSM.scala 1116:48 FSM.scala 1118:33]
  wire [5:0] _GEN_1327 = _T_39 ? 6'hf : _GEN_1317; // @[FSM.scala 1116:48 FSM.scala 1119:35]
  wire [11:0] _GEN_1328 = _T_39 ? {{1'd0}, PEArray_ctrl_2_mask[11:1]} : _GEN_1318; // @[FSM.scala 1116:48 FSM.scala 1120:32]
  wire [7:0] _GEN_1329 = _T_39 ? 8'h40 : _GEN_1319; // @[FSM.scala 1116:48 FSM.scala 1121:41]
  wire [11:0] _GEN_1330 = _T_40 ? 12'h0 : _GEN_1297; // @[FSM.scala 1123:29 FSM.scala 1125:34]
  wire [11:0] _GEN_1331 = _T_40 ? 12'h0 : _GEN_1298; // @[FSM.scala 1123:29 FSM.scala 1125:34]
  wire [11:0] _GEN_1332 = _T_40 ? 12'h0 : _GEN_1328; // @[FSM.scala 1123:29 FSM.scala 1125:34]
  wire [11:0] _GEN_1333 = _T_5 ? _L1_rd_addr_0_T_1 : _GEN_1299; // @[FSM.scala 1130:28 FSM.scala 1132:27]
  wire [11:0] _GEN_1334 = _T_48 ? _L1_rd_addr_0_T_1 : _GEN_1333; // @[FSM.scala 1135:28 FSM.scala 1137:27]
  wire [11:0] _GEN_1335 = _T_48 ? _L1_rd_addr_1_T_1 : _GEN_1300; // @[FSM.scala 1135:28 FSM.scala 1137:27]
  wire [11:0] _GEN_1336 = _T_49 ? _L1_rd_addr_0_T_1 : _GEN_1334; // @[FSM.scala 1140:28 FSM.scala 1142:27]
  wire [11:0] _GEN_1337 = _T_49 ? _L1_rd_addr_1_T_1 : _GEN_1335; // @[FSM.scala 1140:28 FSM.scala 1142:27]
  wire [11:0] _GEN_1338 = _T_49 ? _L1_rd_addr_2_T_1 : _GEN_1301; // @[FSM.scala 1140:28 FSM.scala 1142:27]
  wire [11:0] _GEN_1339 = _T_21 ? _L1_rd_addr_0_T_1 : _GEN_1336; // @[FSM.scala 1145:28 FSM.scala 1147:27]
  wire [11:0] _GEN_1340 = _T_21 ? _L1_rd_addr_1_T_1 : _GEN_1337; // @[FSM.scala 1145:28 FSM.scala 1147:27]
  wire [11:0] _GEN_1341 = _T_21 ? _L1_rd_addr_2_T_1 : _GEN_1338; // @[FSM.scala 1145:28 FSM.scala 1147:27]
  wire [11:0] _GEN_1342 = _T_21 ? _L1_rd_addr_3_T_1 : _GEN_1302; // @[FSM.scala 1145:28 FSM.scala 1147:27]
  wire [11:0] _GEN_1343 = _T_51 ? _L1_rd_addr_0_T_1 : _GEN_1339; // @[FSM.scala 1150:28 FSM.scala 1152:27]
  wire [11:0] _GEN_1344 = _T_51 ? _L1_rd_addr_1_T_1 : _GEN_1340; // @[FSM.scala 1150:28 FSM.scala 1152:27]
  wire [11:0] _GEN_1345 = _T_51 ? _L1_rd_addr_2_T_1 : _GEN_1341; // @[FSM.scala 1150:28 FSM.scala 1152:27]
  wire [11:0] _GEN_1346 = _T_51 ? _L1_rd_addr_3_T_1 : _GEN_1342; // @[FSM.scala 1150:28 FSM.scala 1152:27]
  wire [11:0] _GEN_1347 = _T_51 ? _L1_rd_addr_4_T_1 : _GEN_1303; // @[FSM.scala 1150:28 FSM.scala 1152:27]
  wire [11:0] _GEN_1348 = _T_52 ? _L1_rd_addr_0_T_1 : _GEN_1343; // @[FSM.scala 1155:28 FSM.scala 1157:27]
  wire [11:0] _GEN_1349 = _T_52 ? _L1_rd_addr_1_T_1 : _GEN_1344; // @[FSM.scala 1155:28 FSM.scala 1157:27]
  wire [11:0] _GEN_1350 = _T_52 ? _L1_rd_addr_2_T_1 : _GEN_1345; // @[FSM.scala 1155:28 FSM.scala 1157:27]
  wire [11:0] _GEN_1351 = _T_52 ? _L1_rd_addr_3_T_1 : _GEN_1346; // @[FSM.scala 1155:28 FSM.scala 1157:27]
  wire [11:0] _GEN_1352 = _T_52 ? _L1_rd_addr_4_T_1 : _GEN_1347; // @[FSM.scala 1155:28 FSM.scala 1157:27]
  wire [11:0] _GEN_1353 = _T_52 ? _L1_rd_addr_5_T_1 : _GEN_1304; // @[FSM.scala 1155:28 FSM.scala 1157:27]
  wire [11:0] _GEN_1354 = _T_53 ? _L1_rd_addr_0_T_1 : _GEN_1348; // @[FSM.scala 1160:28 FSM.scala 1162:27]
  wire [11:0] _GEN_1355 = _T_53 ? _L1_rd_addr_1_T_1 : _GEN_1349; // @[FSM.scala 1160:28 FSM.scala 1162:27]
  wire [11:0] _GEN_1356 = _T_53 ? _L1_rd_addr_2_T_1 : _GEN_1350; // @[FSM.scala 1160:28 FSM.scala 1162:27]
  wire [11:0] _GEN_1357 = _T_53 ? _L1_rd_addr_3_T_1 : _GEN_1351; // @[FSM.scala 1160:28 FSM.scala 1162:27]
  wire [11:0] _GEN_1358 = _T_53 ? _L1_rd_addr_4_T_1 : _GEN_1352; // @[FSM.scala 1160:28 FSM.scala 1162:27]
  wire [11:0] _GEN_1359 = _T_53 ? _L1_rd_addr_5_T_1 : _GEN_1353; // @[FSM.scala 1160:28 FSM.scala 1162:27]
  wire [11:0] _GEN_1360 = _T_53 ? _L1_rd_addr_6_T_1 : _GEN_1305; // @[FSM.scala 1160:28 FSM.scala 1162:27]
  wire [11:0] _GEN_1361 = _T_54 ? _L1_rd_addr_0_T_1 : _GEN_1354; // @[FSM.scala 1165:28 FSM.scala 1167:27]
  wire [11:0] _GEN_1362 = _T_54 ? _L1_rd_addr_1_T_1 : _GEN_1355; // @[FSM.scala 1165:28 FSM.scala 1167:27]
  wire [11:0] _GEN_1363 = _T_54 ? _L1_rd_addr_2_T_1 : _GEN_1356; // @[FSM.scala 1165:28 FSM.scala 1167:27]
  wire [11:0] _GEN_1364 = _T_54 ? _L1_rd_addr_3_T_1 : _GEN_1357; // @[FSM.scala 1165:28 FSM.scala 1167:27]
  wire [11:0] _GEN_1365 = _T_54 ? _L1_rd_addr_4_T_1 : _GEN_1358; // @[FSM.scala 1165:28 FSM.scala 1167:27]
  wire [11:0] _GEN_1366 = _T_54 ? _L1_rd_addr_5_T_1 : _GEN_1359; // @[FSM.scala 1165:28 FSM.scala 1167:27]
  wire [11:0] _GEN_1367 = _T_54 ? _L1_rd_addr_6_T_1 : _GEN_1360; // @[FSM.scala 1165:28 FSM.scala 1167:27]
  wire [11:0] _GEN_1368 = _T_54 ? _L1_rd_addr_7_T_1 : _GEN_1306; // @[FSM.scala 1165:28 FSM.scala 1167:27]
  wire [11:0] _GEN_1369 = _T_55 ? _L1_rd_addr_0_T_1 : _GEN_1361; // @[FSM.scala 1170:28 FSM.scala 1172:27]
  wire [11:0] _GEN_1370 = _T_55 ? _L1_rd_addr_1_T_1 : _GEN_1362; // @[FSM.scala 1170:28 FSM.scala 1172:27]
  wire [11:0] _GEN_1371 = _T_55 ? _L1_rd_addr_2_T_1 : _GEN_1363; // @[FSM.scala 1170:28 FSM.scala 1172:27]
  wire [11:0] _GEN_1372 = _T_55 ? _L1_rd_addr_3_T_1 : _GEN_1364; // @[FSM.scala 1170:28 FSM.scala 1172:27]
  wire [11:0] _GEN_1373 = _T_55 ? _L1_rd_addr_4_T_1 : _GEN_1365; // @[FSM.scala 1170:28 FSM.scala 1172:27]
  wire [11:0] _GEN_1374 = _T_55 ? _L1_rd_addr_5_T_1 : _GEN_1366; // @[FSM.scala 1170:28 FSM.scala 1172:27]
  wire [11:0] _GEN_1375 = _T_55 ? _L1_rd_addr_6_T_1 : _GEN_1367; // @[FSM.scala 1170:28 FSM.scala 1172:27]
  wire [11:0] _GEN_1376 = _T_55 ? _L1_rd_addr_7_T_1 : _GEN_1368; // @[FSM.scala 1170:28 FSM.scala 1172:27]
  wire [11:0] _GEN_1377 = _T_55 ? _L1_rd_addr_8_T_1 : _GEN_1307; // @[FSM.scala 1170:28 FSM.scala 1172:27]
  wire [11:0] _GEN_1378 = _T_56 ? _L1_rd_addr_0_T_1 : _GEN_1369; // @[FSM.scala 1175:29 FSM.scala 1177:27]
  wire [11:0] _GEN_1379 = _T_56 ? _L1_rd_addr_1_T_1 : _GEN_1370; // @[FSM.scala 1175:29 FSM.scala 1177:27]
  wire [11:0] _GEN_1380 = _T_56 ? _L1_rd_addr_2_T_1 : _GEN_1371; // @[FSM.scala 1175:29 FSM.scala 1177:27]
  wire [11:0] _GEN_1381 = _T_56 ? _L1_rd_addr_3_T_1 : _GEN_1372; // @[FSM.scala 1175:29 FSM.scala 1177:27]
  wire [11:0] _GEN_1382 = _T_56 ? _L1_rd_addr_4_T_1 : _GEN_1373; // @[FSM.scala 1175:29 FSM.scala 1177:27]
  wire [11:0] _GEN_1383 = _T_56 ? _L1_rd_addr_5_T_1 : _GEN_1374; // @[FSM.scala 1175:29 FSM.scala 1177:27]
  wire [11:0] _GEN_1384 = _T_56 ? _L1_rd_addr_6_T_1 : _GEN_1375; // @[FSM.scala 1175:29 FSM.scala 1177:27]
  wire [11:0] _GEN_1385 = _T_56 ? _L1_rd_addr_7_T_1 : _GEN_1376; // @[FSM.scala 1175:29 FSM.scala 1177:27]
  wire [11:0] _GEN_1386 = _T_56 ? _L1_rd_addr_8_T_1 : _GEN_1377; // @[FSM.scala 1175:29 FSM.scala 1177:27]
  wire [11:0] _GEN_1387 = _T_56 ? _L1_rd_addr_9_T_1 : _GEN_1308; // @[FSM.scala 1175:29 FSM.scala 1177:27]
  wire [11:0] _GEN_1388 = _T_57 ? _L1_rd_addr_0_T_1 : _GEN_1378; // @[FSM.scala 1180:29 FSM.scala 1182:27]
  wire [11:0] _GEN_1389 = _T_57 ? _L1_rd_addr_1_T_1 : _GEN_1379; // @[FSM.scala 1180:29 FSM.scala 1182:27]
  wire [11:0] _GEN_1390 = _T_57 ? _L1_rd_addr_2_T_1 : _GEN_1380; // @[FSM.scala 1180:29 FSM.scala 1182:27]
  wire [11:0] _GEN_1391 = _T_57 ? _L1_rd_addr_3_T_1 : _GEN_1381; // @[FSM.scala 1180:29 FSM.scala 1182:27]
  wire [11:0] _GEN_1392 = _T_57 ? _L1_rd_addr_4_T_1 : _GEN_1382; // @[FSM.scala 1180:29 FSM.scala 1182:27]
  wire [11:0] _GEN_1393 = _T_57 ? _L1_rd_addr_5_T_1 : _GEN_1383; // @[FSM.scala 1180:29 FSM.scala 1182:27]
  wire [11:0] _GEN_1394 = _T_57 ? _L1_rd_addr_6_T_1 : _GEN_1384; // @[FSM.scala 1180:29 FSM.scala 1182:27]
  wire [11:0] _GEN_1395 = _T_57 ? _L1_rd_addr_7_T_1 : _GEN_1385; // @[FSM.scala 1180:29 FSM.scala 1182:27]
  wire [11:0] _GEN_1396 = _T_57 ? _L1_rd_addr_8_T_1 : _GEN_1386; // @[FSM.scala 1180:29 FSM.scala 1182:27]
  wire [11:0] _GEN_1397 = _T_57 ? _L1_rd_addr_9_T_1 : _GEN_1387; // @[FSM.scala 1180:29 FSM.scala 1182:27]
  wire [11:0] _GEN_1398 = _T_57 ? _L1_rd_addr_10_T_1 : _GEN_1309; // @[FSM.scala 1180:29 FSM.scala 1182:27]
  wire  _T_226 = _T_110 & count <= 10'h17f; // @[FSM.scala 1185:30]
  wire [11:0] _GEN_1399 = _T_110 & count <= 10'h17f ? _L1_rd_addr_0_T_1 : _GEN_1388; // @[FSM.scala 1185:50 FSM.scala 1187:27]
  wire [11:0] _GEN_1400 = _T_110 & count <= 10'h17f ? _L1_rd_addr_1_T_1 : _GEN_1389; // @[FSM.scala 1185:50 FSM.scala 1187:27]
  wire [11:0] _GEN_1401 = _T_110 & count <= 10'h17f ? _L1_rd_addr_2_T_1 : _GEN_1390; // @[FSM.scala 1185:50 FSM.scala 1187:27]
  wire [11:0] _GEN_1402 = _T_110 & count <= 10'h17f ? _L1_rd_addr_3_T_1 : _GEN_1391; // @[FSM.scala 1185:50 FSM.scala 1187:27]
  wire [11:0] _GEN_1403 = _T_110 & count <= 10'h17f ? _L1_rd_addr_4_T_1 : _GEN_1392; // @[FSM.scala 1185:50 FSM.scala 1187:27]
  wire [11:0] _GEN_1404 = _T_110 & count <= 10'h17f ? _L1_rd_addr_5_T_1 : _GEN_1393; // @[FSM.scala 1185:50 FSM.scala 1187:27]
  wire [11:0] _GEN_1405 = _T_110 & count <= 10'h17f ? _L1_rd_addr_6_T_1 : _GEN_1394; // @[FSM.scala 1185:50 FSM.scala 1187:27]
  wire [11:0] _GEN_1406 = _T_110 & count <= 10'h17f ? _L1_rd_addr_7_T_1 : _GEN_1395; // @[FSM.scala 1185:50 FSM.scala 1187:27]
  wire [11:0] _GEN_1407 = _T_110 & count <= 10'h17f ? _L1_rd_addr_8_T_1 : _GEN_1396; // @[FSM.scala 1185:50 FSM.scala 1187:27]
  wire [11:0] _GEN_1408 = _T_110 & count <= 10'h17f ? _L1_rd_addr_9_T_1 : _GEN_1397; // @[FSM.scala 1185:50 FSM.scala 1187:27]
  wire [11:0] _GEN_1409 = _T_110 & count <= 10'h17f ? _L1_rd_addr_10_T_1 : _GEN_1398; // @[FSM.scala 1185:50 FSM.scala 1187:27]
  wire [11:0] _GEN_1410 = _T_110 & count <= 10'h17f ? _L1_rd_addr_11_T_1 : _GEN_1310; // @[FSM.scala 1185:50 FSM.scala 1187:27]
  wire  _T_227 = count == 10'h180; // @[FSM.scala 1190:20]
  wire [11:0] _GEN_1411 = count == 10'h180 ? _L1_rd_addr_1_T_1 : _GEN_1400; // @[FSM.scala 1190:30 FSM.scala 1192:27]
  wire [11:0] _GEN_1412 = count == 10'h180 ? _L1_rd_addr_2_T_1 : _GEN_1401; // @[FSM.scala 1190:30 FSM.scala 1192:27]
  wire [11:0] _GEN_1413 = count == 10'h180 ? _L1_rd_addr_3_T_1 : _GEN_1402; // @[FSM.scala 1190:30 FSM.scala 1192:27]
  wire [11:0] _GEN_1414 = count == 10'h180 ? _L1_rd_addr_4_T_1 : _GEN_1403; // @[FSM.scala 1190:30 FSM.scala 1192:27]
  wire [11:0] _GEN_1415 = count == 10'h180 ? _L1_rd_addr_5_T_1 : _GEN_1404; // @[FSM.scala 1190:30 FSM.scala 1192:27]
  wire [11:0] _GEN_1416 = count == 10'h180 ? _L1_rd_addr_6_T_1 : _GEN_1405; // @[FSM.scala 1190:30 FSM.scala 1192:27]
  wire [11:0] _GEN_1417 = count == 10'h180 ? _L1_rd_addr_7_T_1 : _GEN_1406; // @[FSM.scala 1190:30 FSM.scala 1192:27]
  wire [11:0] _GEN_1418 = count == 10'h180 ? _L1_rd_addr_8_T_1 : _GEN_1407; // @[FSM.scala 1190:30 FSM.scala 1192:27]
  wire [11:0] _GEN_1419 = count == 10'h180 ? _L1_rd_addr_9_T_1 : _GEN_1408; // @[FSM.scala 1190:30 FSM.scala 1192:27]
  wire [11:0] _GEN_1420 = count == 10'h180 ? _L1_rd_addr_10_T_1 : _GEN_1409; // @[FSM.scala 1190:30 FSM.scala 1192:27]
  wire [11:0] _GEN_1421 = count == 10'h180 ? _L1_rd_addr_11_T_1 : _GEN_1410; // @[FSM.scala 1190:30 FSM.scala 1192:27]
  wire  _T_228 = count == 10'h181; // @[FSM.scala 1195:20]
  wire [11:0] _GEN_1422 = count == 10'h181 ? _L1_rd_addr_2_T_1 : _GEN_1412; // @[FSM.scala 1195:30 FSM.scala 1197:27]
  wire [11:0] _GEN_1423 = count == 10'h181 ? _L1_rd_addr_3_T_1 : _GEN_1413; // @[FSM.scala 1195:30 FSM.scala 1197:27]
  wire [11:0] _GEN_1424 = count == 10'h181 ? _L1_rd_addr_4_T_1 : _GEN_1414; // @[FSM.scala 1195:30 FSM.scala 1197:27]
  wire [11:0] _GEN_1425 = count == 10'h181 ? _L1_rd_addr_5_T_1 : _GEN_1415; // @[FSM.scala 1195:30 FSM.scala 1197:27]
  wire [11:0] _GEN_1426 = count == 10'h181 ? _L1_rd_addr_6_T_1 : _GEN_1416; // @[FSM.scala 1195:30 FSM.scala 1197:27]
  wire [11:0] _GEN_1427 = count == 10'h181 ? _L1_rd_addr_7_T_1 : _GEN_1417; // @[FSM.scala 1195:30 FSM.scala 1197:27]
  wire [11:0] _GEN_1428 = count == 10'h181 ? _L1_rd_addr_8_T_1 : _GEN_1418; // @[FSM.scala 1195:30 FSM.scala 1197:27]
  wire [11:0] _GEN_1429 = count == 10'h181 ? _L1_rd_addr_9_T_1 : _GEN_1419; // @[FSM.scala 1195:30 FSM.scala 1197:27]
  wire [11:0] _GEN_1430 = count == 10'h181 ? _L1_rd_addr_10_T_1 : _GEN_1420; // @[FSM.scala 1195:30 FSM.scala 1197:27]
  wire [11:0] _GEN_1431 = count == 10'h181 ? _L1_rd_addr_11_T_1 : _GEN_1421; // @[FSM.scala 1195:30 FSM.scala 1197:27]
  wire  _T_229 = count == 10'h182; // @[FSM.scala 1200:20]
  wire [11:0] _GEN_1432 = count == 10'h182 ? _L1_rd_addr_3_T_1 : _GEN_1423; // @[FSM.scala 1200:30 FSM.scala 1202:27]
  wire [11:0] _GEN_1433 = count == 10'h182 ? _L1_rd_addr_4_T_1 : _GEN_1424; // @[FSM.scala 1200:30 FSM.scala 1202:27]
  wire [11:0] _GEN_1434 = count == 10'h182 ? _L1_rd_addr_5_T_1 : _GEN_1425; // @[FSM.scala 1200:30 FSM.scala 1202:27]
  wire [11:0] _GEN_1435 = count == 10'h182 ? _L1_rd_addr_6_T_1 : _GEN_1426; // @[FSM.scala 1200:30 FSM.scala 1202:27]
  wire [11:0] _GEN_1436 = count == 10'h182 ? _L1_rd_addr_7_T_1 : _GEN_1427; // @[FSM.scala 1200:30 FSM.scala 1202:27]
  wire [11:0] _GEN_1437 = count == 10'h182 ? _L1_rd_addr_8_T_1 : _GEN_1428; // @[FSM.scala 1200:30 FSM.scala 1202:27]
  wire [11:0] _GEN_1438 = count == 10'h182 ? _L1_rd_addr_9_T_1 : _GEN_1429; // @[FSM.scala 1200:30 FSM.scala 1202:27]
  wire [11:0] _GEN_1439 = count == 10'h182 ? _L1_rd_addr_10_T_1 : _GEN_1430; // @[FSM.scala 1200:30 FSM.scala 1202:27]
  wire [11:0] _GEN_1440 = count == 10'h182 ? _L1_rd_addr_11_T_1 : _GEN_1431; // @[FSM.scala 1200:30 FSM.scala 1202:27]
  wire  _T_230 = count == 10'h183; // @[FSM.scala 1205:20]
  wire [11:0] _GEN_1441 = count == 10'h183 ? _L1_rd_addr_4_T_1 : _GEN_1433; // @[FSM.scala 1205:30 FSM.scala 1207:27]
  wire [11:0] _GEN_1442 = count == 10'h183 ? _L1_rd_addr_5_T_1 : _GEN_1434; // @[FSM.scala 1205:30 FSM.scala 1207:27]
  wire [11:0] _GEN_1443 = count == 10'h183 ? _L1_rd_addr_6_T_1 : _GEN_1435; // @[FSM.scala 1205:30 FSM.scala 1207:27]
  wire [11:0] _GEN_1444 = count == 10'h183 ? _L1_rd_addr_7_T_1 : _GEN_1436; // @[FSM.scala 1205:30 FSM.scala 1207:27]
  wire [11:0] _GEN_1445 = count == 10'h183 ? _L1_rd_addr_8_T_1 : _GEN_1437; // @[FSM.scala 1205:30 FSM.scala 1207:27]
  wire [11:0] _GEN_1446 = count == 10'h183 ? _L1_rd_addr_9_T_1 : _GEN_1438; // @[FSM.scala 1205:30 FSM.scala 1207:27]
  wire [11:0] _GEN_1447 = count == 10'h183 ? _L1_rd_addr_10_T_1 : _GEN_1439; // @[FSM.scala 1205:30 FSM.scala 1207:27]
  wire [11:0] _GEN_1448 = count == 10'h183 ? _L1_rd_addr_11_T_1 : _GEN_1440; // @[FSM.scala 1205:30 FSM.scala 1207:27]
  wire  _T_231 = count == 10'h184; // @[FSM.scala 1210:20]
  wire [11:0] _GEN_1449 = count == 10'h184 ? _L1_rd_addr_5_T_1 : _GEN_1442; // @[FSM.scala 1210:30 FSM.scala 1212:27]
  wire [11:0] _GEN_1450 = count == 10'h184 ? _L1_rd_addr_6_T_1 : _GEN_1443; // @[FSM.scala 1210:30 FSM.scala 1212:27]
  wire [11:0] _GEN_1451 = count == 10'h184 ? _L1_rd_addr_7_T_1 : _GEN_1444; // @[FSM.scala 1210:30 FSM.scala 1212:27]
  wire [11:0] _GEN_1452 = count == 10'h184 ? _L1_rd_addr_8_T_1 : _GEN_1445; // @[FSM.scala 1210:30 FSM.scala 1212:27]
  wire [11:0] _GEN_1453 = count == 10'h184 ? _L1_rd_addr_9_T_1 : _GEN_1446; // @[FSM.scala 1210:30 FSM.scala 1212:27]
  wire [11:0] _GEN_1454 = count == 10'h184 ? _L1_rd_addr_10_T_1 : _GEN_1447; // @[FSM.scala 1210:30 FSM.scala 1212:27]
  wire [11:0] _GEN_1455 = count == 10'h184 ? _L1_rd_addr_11_T_1 : _GEN_1448; // @[FSM.scala 1210:30 FSM.scala 1212:27]
  wire  _T_232 = count == 10'h185; // @[FSM.scala 1215:20]
  wire [11:0] _GEN_1456 = count == 10'h185 ? _L1_rd_addr_6_T_1 : _GEN_1450; // @[FSM.scala 1215:30 FSM.scala 1217:27]
  wire [11:0] _GEN_1457 = count == 10'h185 ? _L1_rd_addr_7_T_1 : _GEN_1451; // @[FSM.scala 1215:30 FSM.scala 1217:27]
  wire [11:0] _GEN_1458 = count == 10'h185 ? _L1_rd_addr_8_T_1 : _GEN_1452; // @[FSM.scala 1215:30 FSM.scala 1217:27]
  wire [11:0] _GEN_1459 = count == 10'h185 ? _L1_rd_addr_9_T_1 : _GEN_1453; // @[FSM.scala 1215:30 FSM.scala 1217:27]
  wire [11:0] _GEN_1460 = count == 10'h185 ? _L1_rd_addr_10_T_1 : _GEN_1454; // @[FSM.scala 1215:30 FSM.scala 1217:27]
  wire [11:0] _GEN_1461 = count == 10'h185 ? _L1_rd_addr_11_T_1 : _GEN_1455; // @[FSM.scala 1215:30 FSM.scala 1217:27]
  wire  _T_233 = count == 10'h186; // @[FSM.scala 1220:20]
  wire [11:0] _GEN_1462 = count == 10'h186 ? _L1_rd_addr_7_T_1 : _GEN_1457; // @[FSM.scala 1220:30 FSM.scala 1222:27]
  wire [11:0] _GEN_1463 = count == 10'h186 ? _L1_rd_addr_8_T_1 : _GEN_1458; // @[FSM.scala 1220:30 FSM.scala 1222:27]
  wire [11:0] _GEN_1464 = count == 10'h186 ? _L1_rd_addr_9_T_1 : _GEN_1459; // @[FSM.scala 1220:30 FSM.scala 1222:27]
  wire [11:0] _GEN_1465 = count == 10'h186 ? _L1_rd_addr_10_T_1 : _GEN_1460; // @[FSM.scala 1220:30 FSM.scala 1222:27]
  wire [11:0] _GEN_1466 = count == 10'h186 ? _L1_rd_addr_11_T_1 : _GEN_1461; // @[FSM.scala 1220:30 FSM.scala 1222:27]
  wire  _T_234 = count == 10'h187; // @[FSM.scala 1225:20]
  wire [11:0] _GEN_1467 = count == 10'h187 ? _L1_rd_addr_8_T_1 : _GEN_1463; // @[FSM.scala 1225:30 FSM.scala 1227:27]
  wire [11:0] _GEN_1468 = count == 10'h187 ? _L1_rd_addr_9_T_1 : _GEN_1464; // @[FSM.scala 1225:30 FSM.scala 1227:27]
  wire [11:0] _GEN_1469 = count == 10'h187 ? _L1_rd_addr_10_T_1 : _GEN_1465; // @[FSM.scala 1225:30 FSM.scala 1227:27]
  wire [11:0] _GEN_1470 = count == 10'h187 ? _L1_rd_addr_11_T_1 : _GEN_1466; // @[FSM.scala 1225:30 FSM.scala 1227:27]
  wire  _T_235 = count == 10'h188; // @[FSM.scala 1230:20]
  wire [11:0] _GEN_1471 = count == 10'h188 ? _L1_rd_addr_9_T_1 : _GEN_1468; // @[FSM.scala 1230:30 FSM.scala 1232:27]
  wire [11:0] _GEN_1472 = count == 10'h188 ? _L1_rd_addr_10_T_1 : _GEN_1469; // @[FSM.scala 1230:30 FSM.scala 1232:27]
  wire [11:0] _GEN_1473 = count == 10'h188 ? _L1_rd_addr_11_T_1 : _GEN_1470; // @[FSM.scala 1230:30 FSM.scala 1232:27]
  wire  _T_236 = count == 10'h189; // @[FSM.scala 1235:20]
  wire [11:0] _GEN_1474 = count == 10'h189 ? _L1_rd_addr_10_T_1 : _GEN_1472; // @[FSM.scala 1235:30 FSM.scala 1237:27]
  wire [11:0] _GEN_1475 = count == 10'h189 ? _L1_rd_addr_11_T_1 : _GEN_1473; // @[FSM.scala 1235:30 FSM.scala 1237:27]
  wire [11:0] _GEN_1476 = _T_65 ? _L1_rd_addr_11_T_1 : _GEN_1475; // @[FSM.scala 1240:30 FSM.scala 1242:27]
  wire  _T_240 = _T_124 & count <= 10'h18d; // @[FSM.scala 1246:30]
  wire [5:0] _Uhht_1_wrAddr_T_1 = Uhht_1_wrAddr + 6'h1; // @[FSM.scala 1252:46]
  wire [5:0] _GEN_1477 = _T_127 ? 6'h0 : _Uhht_1_wrAddr_T_1; // @[FSM.scala 1247:33 FSM.scala 1248:27 FSM.scala 1252:29]
  wire [5:0] _GEN_1479 = _T_124 & count <= 10'h18d ? _GEN_1477 : _GEN_1322; // @[FSM.scala 1246:50]
  wire  _GEN_1480 = _T_124 & count <= 10'h18d | Uhht_1_wrEna; // @[FSM.scala 1246:50 FSM.scala 91:36]
  wire [9:0] _GEN_1481 = _T_69 ? 10'h0 : _GEN_1313; // @[FSM.scala 1257:30 FSM.scala 1258:17]
  wire [6:0] _GEN_1482 = _T_69 ? 7'h0 : _GEN_702; // @[FSM.scala 1257:30 FSM.scala 1259:18]
  wire  _GEN_1483 = _T_69 ? 1'h0 : _GEN_1480; // @[FSM.scala 1257:30 FSM.scala 1260:24]
  wire [3:0] _GEN_1484 = _T_69 ? 4'h5 : _GEN_1312; // @[FSM.scala 1257:30 FSM.scala 1261:21]
  wire [9:0] _GEN_1485 = gru_state == 4'h4 ? _GEN_1481 : _GEN_1285; // @[FSM.scala 1085:30]
  wire [6:0] _GEN_1486 = gru_state == 4'h4 ? _GEN_1482 : _GEN_1286; // @[FSM.scala 1085:30]
  wire [2:0] _GEN_1487 = gru_state == 4'h4 ? _GEN_1325 : _GEN_1287; // @[FSM.scala 1085:30]
  wire [9:0] _GEN_1488 = gru_state == 4'h4 ? _GEN_1326 : _GEN_1288; // @[FSM.scala 1085:30]
  wire [5:0] _GEN_1489 = gru_state == 4'h4 ? _GEN_1327 : _GEN_1289; // @[FSM.scala 1085:30]
  wire [11:0] _GEN_1490 = gru_state == 4'h4 ? _GEN_1332 : _GEN_1290; // @[FSM.scala 1085:30]
  wire [7:0] _GEN_1491 = gru_state == 4'h4 ? _GEN_1329 : _GEN_1291; // @[FSM.scala 1085:30]
  wire [1:0] _GEN_1492 = gru_state == 4'h4 ? _GEN_1320 : _GEN_1292; // @[FSM.scala 1085:30]
  wire [3:0] _GEN_1493 = gru_state == 4'h4 ? _GEN_1321 : _GEN_1293; // @[FSM.scala 1085:30]
  wire [5:0] _GEN_1494 = gru_state == 4'h4 ? _GEN_1479 : Uhht_1_wrAddr; // @[FSM.scala 1085:30 FSM.scala 92:36]
  wire [1:0] _GEN_1495 = gru_state == 4'h4 ? _GEN_1323 : _GEN_1295; // @[FSM.scala 1085:30]
  wire [1:0] _GEN_1496 = gru_state == 4'h4 ? _GEN_1324 : _GEN_1296; // @[FSM.scala 1085:30]
  wire [11:0] _GEN_1497 = gru_state == 4'h4 ? _GEN_1330 : _GEN_1297; // @[FSM.scala 1085:30]
  wire [11:0] _GEN_1498 = gru_state == 4'h4 ? _GEN_1331 : _GEN_1298; // @[FSM.scala 1085:30]
  wire [11:0] _GEN_1499 = gru_state == 4'h4 ? _GEN_1399 : _GEN_1299; // @[FSM.scala 1085:30]
  wire [11:0] _GEN_1500 = gru_state == 4'h4 ? _GEN_1411 : _GEN_1300; // @[FSM.scala 1085:30]
  wire [11:0] _GEN_1501 = gru_state == 4'h4 ? _GEN_1422 : _GEN_1301; // @[FSM.scala 1085:30]
  wire [11:0] _GEN_1502 = gru_state == 4'h4 ? _GEN_1432 : _GEN_1302; // @[FSM.scala 1085:30]
  wire [11:0] _GEN_1503 = gru_state == 4'h4 ? _GEN_1441 : _GEN_1303; // @[FSM.scala 1085:30]
  wire [11:0] _GEN_1504 = gru_state == 4'h4 ? _GEN_1449 : _GEN_1304; // @[FSM.scala 1085:30]
  wire [11:0] _GEN_1505 = gru_state == 4'h4 ? _GEN_1456 : _GEN_1305; // @[FSM.scala 1085:30]
  wire [11:0] _GEN_1506 = gru_state == 4'h4 ? _GEN_1462 : _GEN_1306; // @[FSM.scala 1085:30]
  wire [11:0] _GEN_1507 = gru_state == 4'h4 ? _GEN_1467 : _GEN_1307; // @[FSM.scala 1085:30]
  wire [11:0] _GEN_1508 = gru_state == 4'h4 ? _GEN_1471 : _GEN_1308; // @[FSM.scala 1085:30]
  wire [11:0] _GEN_1509 = gru_state == 4'h4 ? _GEN_1474 : _GEN_1309; // @[FSM.scala 1085:30]
  wire [11:0] _GEN_1510 = gru_state == 4'h4 ? _GEN_1476 : _GEN_1310; // @[FSM.scala 1085:30]
  wire  _GEN_1511 = gru_state == 4'h4 ? _GEN_1483 : Uhht_1_wrEna; // @[FSM.scala 1085:30 FSM.scala 91:36]
  wire [3:0] _GEN_1512 = gru_state == 4'h4 ? _GEN_1484 : _GEN_1312; // @[FSM.scala 1085:30]
  wire [9:0] _GEN_1513 = count != 10'h44 ? _count_T_1 : _GEN_1485; // @[FSM.scala 1266:29 FSM.scala 1267:17]
  wire [5:0] _GEN_1514 = _T_3 ? 6'h0 : Zt_rdAddr; // @[FSM.scala 1270:28 FSM.scala 1271:21 FSM.scala 81:36]
  wire [5:0] _GEN_1515 = _T_3 ? 6'h0 : Rt_rdAddr; // @[FSM.scala 1270:28 FSM.scala 1272:21 FSM.scala 84:36]
  wire [5:0] _GEN_1516 = _T_3 ? 6'h0 : WhXt_rdAddr; // @[FSM.scala 1270:28 FSM.scala 1273:23 FSM.scala 87:36]
  wire [5:0] _GEN_1517 = _T_3 ? 6'h0 : Uhht_1_rdAddr; // @[FSM.scala 1270:28 FSM.scala 1274:25 FSM.scala 90:36]
  wire [5:0] _Zt_rdAddr_T_1 = Zt_rdAddr + 6'h1; // @[FSM.scala 1277:34]
  wire [5:0] _Rt_rdAddr_T_1 = Rt_rdAddr + 6'h1; // @[FSM.scala 1278:34]
  wire [5:0] _WhXt_rdAddr_T_1 = WhXt_rdAddr + 6'h1; // @[FSM.scala 1279:38]
  wire [5:0] _Uhht_1_rdAddr_T_1 = Uhht_1_rdAddr + 6'h1; // @[FSM.scala 1280:42]
  wire [5:0] _GEN_1518 = _T_18 & count <= 10'h3f ? _Zt_rdAddr_T_1 : _GEN_1514; // @[FSM.scala 1276:48 FSM.scala 1277:21]
  wire [5:0] _GEN_1519 = _T_18 & count <= 10'h3f ? _Rt_rdAddr_T_1 : _GEN_1515; // @[FSM.scala 1276:48 FSM.scala 1278:21]
  wire [5:0] _GEN_1520 = _T_18 & count <= 10'h3f ? _WhXt_rdAddr_T_1 : _GEN_1516; // @[FSM.scala 1276:48 FSM.scala 1279:23]
  wire [5:0] _GEN_1521 = _T_18 & count <= 10'h3f ? _Uhht_1_rdAddr_T_1 : _GEN_1517; // @[FSM.scala 1276:48 FSM.scala 1280:25]
  wire [5:0] _GEN_1522 = _T_49 ? 6'h0 : Ht_wrAddr; // @[FSM.scala 1283:28 FSM.scala 1284:21 FSM.scala 80:36]
  wire  _GEN_1523 = _T_49 | Ht_wrEna; // @[FSM.scala 1283:28 FSM.scala 1285:20 FSM.scala 79:36]
  wire [5:0] _Ht_wrAddr_T_1 = Ht_wrAddr + 6'h1; // @[FSM.scala 1288:34]
  wire [5:0] _GEN_1524 = count <= 10'h4 & count >= 10'h43 ? _Ht_wrAddr_T_1 : _GEN_1522; // @[FSM.scala 1287:44 FSM.scala 1288:21]
  wire [5:0] _gru_count_T_1 = gru_count + 6'h1; // @[FSM.scala 1299:36]
  wire [2:0] _GEN_1525 = gru_count == 6'h3f ? 3'h5 : 3'h4; // @[FSM.scala 1294:35 FSM.scala 1295:19 FSM.scala 1298:19]
  wire [5:0] _GEN_1526 = gru_count == 6'h3f ? 6'h0 : _gru_count_T_1; // @[FSM.scala 1294:35 FSM.scala 1296:23 FSM.scala 1299:23]
  wire [9:0] _GEN_1527 = count == 10'h44 ? 10'h0 : _GEN_1513; // @[FSM.scala 1290:29 FSM.scala 1291:17]
  wire  _GEN_1528 = count == 10'h44 ? 1'h0 : _GEN_1523; // @[FSM.scala 1290:29 FSM.scala 1292:20]
  wire [3:0] _GEN_1529 = count == 10'h44 ? 4'h0 : _GEN_1512; // @[FSM.scala 1290:29 FSM.scala 1293:21]
  wire [2:0] _GEN_1530 = count == 10'h44 ? _GEN_1525 : state; // @[FSM.scala 1290:29 FSM.scala 159:22]
  wire [5:0] _GEN_1531 = count == 10'h44 ? _GEN_1526 : gru_count; // @[FSM.scala 1290:29 FSM.scala 164:26]
  wire [9:0] _GEN_1532 = gru_state == 4'h5 ? _GEN_1527 : _GEN_1485; // @[FSM.scala 1265:30]
  wire [5:0] _GEN_1533 = gru_state == 4'h5 ? _GEN_1518 : Zt_rdAddr; // @[FSM.scala 1265:30 FSM.scala 81:36]
  wire [5:0] _GEN_1534 = gru_state == 4'h5 ? _GEN_1519 : Rt_rdAddr; // @[FSM.scala 1265:30 FSM.scala 84:36]
  wire [5:0] _GEN_1535 = gru_state == 4'h5 ? _GEN_1520 : WhXt_rdAddr; // @[FSM.scala 1265:30 FSM.scala 87:36]
  wire [5:0] _GEN_1536 = gru_state == 4'h5 ? _GEN_1521 : Uhht_1_rdAddr; // @[FSM.scala 1265:30 FSM.scala 90:36]
  wire [5:0] _GEN_1537 = gru_state == 4'h5 ? _GEN_1524 : Ht_wrAddr; // @[FSM.scala 1265:30 FSM.scala 80:36]
  wire  _GEN_1538 = gru_state == 4'h5 ? _GEN_1528 : Ht_wrEna; // @[FSM.scala 1265:30 FSM.scala 79:36]
  wire [3:0] _GEN_1539 = gru_state == 4'h5 ? _GEN_1529 : _GEN_1512; // @[FSM.scala 1265:30]
  wire [2:0] _GEN_1540 = gru_state == 4'h5 ? _GEN_1530 : state; // @[FSM.scala 1265:30 FSM.scala 159:22]
  wire [5:0] _GEN_1541 = gru_state == 4'h5 ? _GEN_1531 : gru_count; // @[FSM.scala 1265:30 FSM.scala 164:26]
  wire  _T_255 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _T_257 = count != 10'ha; // @[FSM.scala 1307:20]
  wire [9:0] _GEN_1542 = count != 10'ha ? _count_T_1 : count; // @[FSM.scala 1307:29 FSM.scala 1308:17 FSM.scala 161:22]
  wire [9:0] _GEN_1545 = _T_3 ? 10'h7 : PEArray_ctrl_2_count; // @[FSM.scala 1311:28 FSM.scala 1315:33 FSM.scala 64:28]
  wire [9:0] _GEN_1554 = _T_56 ? 10'h0 : _GEN_1542; // @[FSM.scala 1333:29 FSM.scala 1334:17]
  wire [1:0] _GEN_1555 = _T_56 ? 2'h1 : fc_state; // @[FSM.scala 1333:29 FSM.scala 1335:20 FSM.scala 166:25]
  wire [9:0] _GEN_1556 = fc_state == 2'h0 ? _GEN_1554 : count; // @[FSM.scala 1306:29 FSM.scala 161:22]
  wire [2:0] _GEN_1557 = fc_state == 2'h0 ? _GEN_640 : PEArray_ctrl_2_control; // @[FSM.scala 1306:29 FSM.scala 64:28]
  wire [11:0] _GEN_1558 = fc_state == 2'h0 ? _GEN_108 : PEArray_ctrl_2_mask; // @[FSM.scala 1306:29 FSM.scala 64:28]
  wire [9:0] _GEN_1559 = fc_state == 2'h0 ? _GEN_1545 : PEArray_ctrl_2_count; // @[FSM.scala 1306:29 FSM.scala 64:28]
  wire [5:0] _GEN_1560 = fc_state == 2'h0 ? _GEN_643 : PEArray_ctrl_2_L0index; // @[FSM.scala 1306:29 FSM.scala 64:28]
  wire [1:0] _GEN_1561 = fc_state == 2'h0 ? _GEN_644 : PE_above_data_ctrl; // @[FSM.scala 1306:29 FSM.scala 74:35]
  wire [3:0] _GEN_1562 = fc_state == 2'h0 ? _GEN_105 : PE_rd_data_mux; // @[FSM.scala 1306:29 FSM.scala 61:32]
  wire [11:0] _GEN_1563 = fc_state == 2'h0 ? _GEN_646 : PEArray_ctrl_0_mask; // @[FSM.scala 1306:29 FSM.scala 64:28]
  wire [11:0] _GEN_1564 = fc_state == 2'h0 ? _GEN_647 : PEArray_ctrl_1_mask; // @[FSM.scala 1306:29 FSM.scala 64:28]
  wire [2:0] _GEN_1565 = fc_state == 2'h0 ? _GEN_650 : Ht_to_PE_control; // @[FSM.scala 1306:29 FSM.scala 77:36]
  wire [1:0] _GEN_1566 = fc_state == 2'h0 ? _GEN_1555 : fc_state; // @[FSM.scala 1306:29 FSM.scala 166:25]
  wire [9:0] _GEN_1567 = _T_206 ? _count_T_1 : _GEN_1556; // @[FSM.scala 1339:30 FSM.scala 1340:17]
  wire [2:0] _GEN_1569 = _T_3 ? 3'h4 : _GEN_1557; // @[FSM.scala 1350:28 FSM.scala 1352:35]
  wire [9:0] _GEN_1570 = _T_3 ? 10'h17f : _GEN_1559; // @[FSM.scala 1350:28 FSM.scala 1353:33]
  wire [5:0] _GEN_1571 = _T_3 ? 6'hf : _GEN_1560; // @[FSM.scala 1350:28 FSM.scala 1354:35]
  wire [11:0] _GEN_1572 = _T_3 ? 12'h800 : _GEN_1558; // @[FSM.scala 1350:28 FSM.scala 1355:32]
  wire [1:0] _GEN_1574 = _T_3 ? 2'h0 : _GEN_1561; // @[FSM.scala 1350:28 FSM.scala 1359:30]
  wire [3:0] _GEN_1575 = _T_3 ? 4'h0 : _GEN_1562; // @[FSM.scala 1350:28 FSM.scala 1360:26]
  wire [5:0] _GEN_1576 = _T_3 ? 6'h0 : FC_temp_wrAddr; // @[FSM.scala 1350:28 FSM.scala 1363:26 FSM.scala 97:38]
  wire [1:0] _GEN_1577 = _T_3 ? 2'h3 : BN_Unit_ctrl; // @[FSM.scala 1350:28 FSM.scala 1364:24 FSM.scala 69:28]
  wire [1:0] _GEN_1578 = _T_3 ? 2'h3 : Activation_ctrl; // @[FSM.scala 1350:28 FSM.scala 1365:27 FSM.scala 75:32]
  wire [2:0] _GEN_1579 = _T_39 ? 3'h4 : _GEN_1569; // @[FSM.scala 1369:48 FSM.scala 1370:35]
  wire [9:0] _GEN_1580 = _T_39 ? 10'h17f : _GEN_1570; // @[FSM.scala 1369:48 FSM.scala 1371:33]
  wire [5:0] _GEN_1581 = _T_39 ? 6'hf : _GEN_1571; // @[FSM.scala 1369:48 FSM.scala 1372:35]
  wire [11:0] _GEN_1582 = _T_39 ? {{1'd0}, PEArray_ctrl_2_mask[11:1]} : _GEN_1572; // @[FSM.scala 1369:48 FSM.scala 1373:32]
  wire [11:0] _GEN_1584 = _T_40 ? 12'h0 : _GEN_1563; // @[FSM.scala 1376:29 FSM.scala 1378:34]
  wire [11:0] _GEN_1585 = _T_40 ? 12'h0 : _GEN_1564; // @[FSM.scala 1376:29 FSM.scala 1378:34]
  wire [11:0] _GEN_1586 = _T_40 ? 12'h0 : _GEN_1582; // @[FSM.scala 1376:29 FSM.scala 1378:34]
  wire [11:0] _GEN_1587 = _T_5 ? _L1_rd_addr_0_T_1 : L1_rd_addr_0; // @[FSM.scala 1383:28 FSM.scala 1385:27 FSM.scala 60:28]
  wire [11:0] _GEN_1588 = _T_48 ? _L1_rd_addr_0_T_1 : _GEN_1587; // @[FSM.scala 1388:28 FSM.scala 1390:27]
  wire [11:0] _GEN_1589 = _T_48 ? _L1_rd_addr_1_T_1 : L1_rd_addr_1; // @[FSM.scala 1388:28 FSM.scala 1390:27 FSM.scala 60:28]
  wire [11:0] _GEN_1590 = _T_49 ? _L1_rd_addr_0_T_1 : _GEN_1588; // @[FSM.scala 1393:28 FSM.scala 1395:27]
  wire [11:0] _GEN_1591 = _T_49 ? _L1_rd_addr_1_T_1 : _GEN_1589; // @[FSM.scala 1393:28 FSM.scala 1395:27]
  wire [11:0] _GEN_1592 = _T_49 ? _L1_rd_addr_2_T_1 : L1_rd_addr_2; // @[FSM.scala 1393:28 FSM.scala 1395:27 FSM.scala 60:28]
  wire [11:0] _GEN_1593 = _T_21 ? _L1_rd_addr_0_T_1 : _GEN_1590; // @[FSM.scala 1398:28 FSM.scala 1400:27]
  wire [11:0] _GEN_1594 = _T_21 ? _L1_rd_addr_1_T_1 : _GEN_1591; // @[FSM.scala 1398:28 FSM.scala 1400:27]
  wire [11:0] _GEN_1595 = _T_21 ? _L1_rd_addr_2_T_1 : _GEN_1592; // @[FSM.scala 1398:28 FSM.scala 1400:27]
  wire [11:0] _GEN_1596 = _T_21 ? _L1_rd_addr_3_T_1 : L1_rd_addr_3; // @[FSM.scala 1398:28 FSM.scala 1400:27 FSM.scala 60:28]
  wire [11:0] _GEN_1597 = _T_51 ? _L1_rd_addr_0_T_1 : _GEN_1593; // @[FSM.scala 1403:28 FSM.scala 1405:27]
  wire [11:0] _GEN_1598 = _T_51 ? _L1_rd_addr_1_T_1 : _GEN_1594; // @[FSM.scala 1403:28 FSM.scala 1405:27]
  wire [11:0] _GEN_1599 = _T_51 ? _L1_rd_addr_2_T_1 : _GEN_1595; // @[FSM.scala 1403:28 FSM.scala 1405:27]
  wire [11:0] _GEN_1600 = _T_51 ? _L1_rd_addr_3_T_1 : _GEN_1596; // @[FSM.scala 1403:28 FSM.scala 1405:27]
  wire [11:0] _GEN_1601 = _T_51 ? _L1_rd_addr_4_T_1 : L1_rd_addr_4; // @[FSM.scala 1403:28 FSM.scala 1405:27 FSM.scala 60:28]
  wire [11:0] _GEN_1602 = _T_52 ? _L1_rd_addr_0_T_1 : _GEN_1597; // @[FSM.scala 1408:28 FSM.scala 1410:27]
  wire [11:0] _GEN_1603 = _T_52 ? _L1_rd_addr_1_T_1 : _GEN_1598; // @[FSM.scala 1408:28 FSM.scala 1410:27]
  wire [11:0] _GEN_1604 = _T_52 ? _L1_rd_addr_2_T_1 : _GEN_1599; // @[FSM.scala 1408:28 FSM.scala 1410:27]
  wire [11:0] _GEN_1605 = _T_52 ? _L1_rd_addr_3_T_1 : _GEN_1600; // @[FSM.scala 1408:28 FSM.scala 1410:27]
  wire [11:0] _GEN_1606 = _T_52 ? _L1_rd_addr_4_T_1 : _GEN_1601; // @[FSM.scala 1408:28 FSM.scala 1410:27]
  wire [11:0] _GEN_1607 = _T_52 ? _L1_rd_addr_5_T_1 : L1_rd_addr_5; // @[FSM.scala 1408:28 FSM.scala 1410:27 FSM.scala 60:28]
  wire [11:0] _GEN_1608 = _T_53 ? _L1_rd_addr_0_T_1 : _GEN_1602; // @[FSM.scala 1413:28 FSM.scala 1415:27]
  wire [11:0] _GEN_1609 = _T_53 ? _L1_rd_addr_1_T_1 : _GEN_1603; // @[FSM.scala 1413:28 FSM.scala 1415:27]
  wire [11:0] _GEN_1610 = _T_53 ? _L1_rd_addr_2_T_1 : _GEN_1604; // @[FSM.scala 1413:28 FSM.scala 1415:27]
  wire [11:0] _GEN_1611 = _T_53 ? _L1_rd_addr_3_T_1 : _GEN_1605; // @[FSM.scala 1413:28 FSM.scala 1415:27]
  wire [11:0] _GEN_1612 = _T_53 ? _L1_rd_addr_4_T_1 : _GEN_1606; // @[FSM.scala 1413:28 FSM.scala 1415:27]
  wire [11:0] _GEN_1613 = _T_53 ? _L1_rd_addr_5_T_1 : _GEN_1607; // @[FSM.scala 1413:28 FSM.scala 1415:27]
  wire [11:0] _GEN_1614 = _T_53 ? _L1_rd_addr_6_T_1 : L1_rd_addr_6; // @[FSM.scala 1413:28 FSM.scala 1415:27 FSM.scala 60:28]
  wire [11:0] _GEN_1615 = _T_54 ? _L1_rd_addr_0_T_1 : _GEN_1608; // @[FSM.scala 1418:28 FSM.scala 1420:27]
  wire [11:0] _GEN_1616 = _T_54 ? _L1_rd_addr_1_T_1 : _GEN_1609; // @[FSM.scala 1418:28 FSM.scala 1420:27]
  wire [11:0] _GEN_1617 = _T_54 ? _L1_rd_addr_2_T_1 : _GEN_1610; // @[FSM.scala 1418:28 FSM.scala 1420:27]
  wire [11:0] _GEN_1618 = _T_54 ? _L1_rd_addr_3_T_1 : _GEN_1611; // @[FSM.scala 1418:28 FSM.scala 1420:27]
  wire [11:0] _GEN_1619 = _T_54 ? _L1_rd_addr_4_T_1 : _GEN_1612; // @[FSM.scala 1418:28 FSM.scala 1420:27]
  wire [11:0] _GEN_1620 = _T_54 ? _L1_rd_addr_5_T_1 : _GEN_1613; // @[FSM.scala 1418:28 FSM.scala 1420:27]
  wire [11:0] _GEN_1621 = _T_54 ? _L1_rd_addr_6_T_1 : _GEN_1614; // @[FSM.scala 1418:28 FSM.scala 1420:27]
  wire [11:0] _GEN_1622 = _T_54 ? _L1_rd_addr_7_T_1 : L1_rd_addr_7; // @[FSM.scala 1418:28 FSM.scala 1420:27 FSM.scala 60:28]
  wire [11:0] _GEN_1623 = _T_55 ? _L1_rd_addr_0_T_1 : _GEN_1615; // @[FSM.scala 1423:28 FSM.scala 1425:27]
  wire [11:0] _GEN_1624 = _T_55 ? _L1_rd_addr_1_T_1 : _GEN_1616; // @[FSM.scala 1423:28 FSM.scala 1425:27]
  wire [11:0] _GEN_1625 = _T_55 ? _L1_rd_addr_2_T_1 : _GEN_1617; // @[FSM.scala 1423:28 FSM.scala 1425:27]
  wire [11:0] _GEN_1626 = _T_55 ? _L1_rd_addr_3_T_1 : _GEN_1618; // @[FSM.scala 1423:28 FSM.scala 1425:27]
  wire [11:0] _GEN_1627 = _T_55 ? _L1_rd_addr_4_T_1 : _GEN_1619; // @[FSM.scala 1423:28 FSM.scala 1425:27]
  wire [11:0] _GEN_1628 = _T_55 ? _L1_rd_addr_5_T_1 : _GEN_1620; // @[FSM.scala 1423:28 FSM.scala 1425:27]
  wire [11:0] _GEN_1629 = _T_55 ? _L1_rd_addr_6_T_1 : _GEN_1621; // @[FSM.scala 1423:28 FSM.scala 1425:27]
  wire [11:0] _GEN_1630 = _T_55 ? _L1_rd_addr_7_T_1 : _GEN_1622; // @[FSM.scala 1423:28 FSM.scala 1425:27]
  wire [11:0] _GEN_1631 = _T_55 ? _L1_rd_addr_8_T_1 : L1_rd_addr_8; // @[FSM.scala 1423:28 FSM.scala 1425:27 FSM.scala 60:28]
  wire [11:0] _GEN_1632 = _T_56 ? _L1_rd_addr_0_T_1 : _GEN_1623; // @[FSM.scala 1428:29 FSM.scala 1430:27]
  wire [11:0] _GEN_1633 = _T_56 ? _L1_rd_addr_1_T_1 : _GEN_1624; // @[FSM.scala 1428:29 FSM.scala 1430:27]
  wire [11:0] _GEN_1634 = _T_56 ? _L1_rd_addr_2_T_1 : _GEN_1625; // @[FSM.scala 1428:29 FSM.scala 1430:27]
  wire [11:0] _GEN_1635 = _T_56 ? _L1_rd_addr_3_T_1 : _GEN_1626; // @[FSM.scala 1428:29 FSM.scala 1430:27]
  wire [11:0] _GEN_1636 = _T_56 ? _L1_rd_addr_4_T_1 : _GEN_1627; // @[FSM.scala 1428:29 FSM.scala 1430:27]
  wire [11:0] _GEN_1637 = _T_56 ? _L1_rd_addr_5_T_1 : _GEN_1628; // @[FSM.scala 1428:29 FSM.scala 1430:27]
  wire [11:0] _GEN_1638 = _T_56 ? _L1_rd_addr_6_T_1 : _GEN_1629; // @[FSM.scala 1428:29 FSM.scala 1430:27]
  wire [11:0] _GEN_1639 = _T_56 ? _L1_rd_addr_7_T_1 : _GEN_1630; // @[FSM.scala 1428:29 FSM.scala 1430:27]
  wire [11:0] _GEN_1640 = _T_56 ? _L1_rd_addr_8_T_1 : _GEN_1631; // @[FSM.scala 1428:29 FSM.scala 1430:27]
  wire [11:0] _GEN_1641 = _T_56 ? _L1_rd_addr_9_T_1 : L1_rd_addr_9; // @[FSM.scala 1428:29 FSM.scala 1430:27 FSM.scala 60:28]
  wire [11:0] _GEN_1642 = _T_57 ? _L1_rd_addr_0_T_1 : _GEN_1632; // @[FSM.scala 1433:29 FSM.scala 1435:27]
  wire [11:0] _GEN_1643 = _T_57 ? _L1_rd_addr_1_T_1 : _GEN_1633; // @[FSM.scala 1433:29 FSM.scala 1435:27]
  wire [11:0] _GEN_1644 = _T_57 ? _L1_rd_addr_2_T_1 : _GEN_1634; // @[FSM.scala 1433:29 FSM.scala 1435:27]
  wire [11:0] _GEN_1645 = _T_57 ? _L1_rd_addr_3_T_1 : _GEN_1635; // @[FSM.scala 1433:29 FSM.scala 1435:27]
  wire [11:0] _GEN_1646 = _T_57 ? _L1_rd_addr_4_T_1 : _GEN_1636; // @[FSM.scala 1433:29 FSM.scala 1435:27]
  wire [11:0] _GEN_1647 = _T_57 ? _L1_rd_addr_5_T_1 : _GEN_1637; // @[FSM.scala 1433:29 FSM.scala 1435:27]
  wire [11:0] _GEN_1648 = _T_57 ? _L1_rd_addr_6_T_1 : _GEN_1638; // @[FSM.scala 1433:29 FSM.scala 1435:27]
  wire [11:0] _GEN_1649 = _T_57 ? _L1_rd_addr_7_T_1 : _GEN_1639; // @[FSM.scala 1433:29 FSM.scala 1435:27]
  wire [11:0] _GEN_1650 = _T_57 ? _L1_rd_addr_8_T_1 : _GEN_1640; // @[FSM.scala 1433:29 FSM.scala 1435:27]
  wire [11:0] _GEN_1651 = _T_57 ? _L1_rd_addr_9_T_1 : _GEN_1641; // @[FSM.scala 1433:29 FSM.scala 1435:27]
  wire [11:0] _GEN_1652 = _T_57 ? _L1_rd_addr_10_T_1 : L1_rd_addr_10; // @[FSM.scala 1433:29 FSM.scala 1435:27 FSM.scala 60:28]
  wire [11:0] _GEN_1653 = _T_226 ? _L1_rd_addr_0_T_1 : _GEN_1642; // @[FSM.scala 1438:50 FSM.scala 1440:27]
  wire [11:0] _GEN_1654 = _T_226 ? _L1_rd_addr_1_T_1 : _GEN_1643; // @[FSM.scala 1438:50 FSM.scala 1440:27]
  wire [11:0] _GEN_1655 = _T_226 ? _L1_rd_addr_2_T_1 : _GEN_1644; // @[FSM.scala 1438:50 FSM.scala 1440:27]
  wire [11:0] _GEN_1656 = _T_226 ? _L1_rd_addr_3_T_1 : _GEN_1645; // @[FSM.scala 1438:50 FSM.scala 1440:27]
  wire [11:0] _GEN_1657 = _T_226 ? _L1_rd_addr_4_T_1 : _GEN_1646; // @[FSM.scala 1438:50 FSM.scala 1440:27]
  wire [11:0] _GEN_1658 = _T_226 ? _L1_rd_addr_5_T_1 : _GEN_1647; // @[FSM.scala 1438:50 FSM.scala 1440:27]
  wire [11:0] _GEN_1659 = _T_226 ? _L1_rd_addr_6_T_1 : _GEN_1648; // @[FSM.scala 1438:50 FSM.scala 1440:27]
  wire [11:0] _GEN_1660 = _T_226 ? _L1_rd_addr_7_T_1 : _GEN_1649; // @[FSM.scala 1438:50 FSM.scala 1440:27]
  wire [11:0] _GEN_1661 = _T_226 ? _L1_rd_addr_8_T_1 : _GEN_1650; // @[FSM.scala 1438:50 FSM.scala 1440:27]
  wire [11:0] _GEN_1662 = _T_226 ? _L1_rd_addr_9_T_1 : _GEN_1651; // @[FSM.scala 1438:50 FSM.scala 1440:27]
  wire [11:0] _GEN_1663 = _T_226 ? _L1_rd_addr_10_T_1 : _GEN_1652; // @[FSM.scala 1438:50 FSM.scala 1440:27]
  wire [11:0] _GEN_1664 = _T_226 ? _L1_rd_addr_11_T_1 : L1_rd_addr_11; // @[FSM.scala 1438:50 FSM.scala 1440:27 FSM.scala 60:28]
  wire [11:0] _GEN_1665 = _T_227 ? _L1_rd_addr_1_T_1 : _GEN_1654; // @[FSM.scala 1443:30 FSM.scala 1445:27]
  wire [11:0] _GEN_1666 = _T_227 ? _L1_rd_addr_2_T_1 : _GEN_1655; // @[FSM.scala 1443:30 FSM.scala 1445:27]
  wire [11:0] _GEN_1667 = _T_227 ? _L1_rd_addr_3_T_1 : _GEN_1656; // @[FSM.scala 1443:30 FSM.scala 1445:27]
  wire [11:0] _GEN_1668 = _T_227 ? _L1_rd_addr_4_T_1 : _GEN_1657; // @[FSM.scala 1443:30 FSM.scala 1445:27]
  wire [11:0] _GEN_1669 = _T_227 ? _L1_rd_addr_5_T_1 : _GEN_1658; // @[FSM.scala 1443:30 FSM.scala 1445:27]
  wire [11:0] _GEN_1670 = _T_227 ? _L1_rd_addr_6_T_1 : _GEN_1659; // @[FSM.scala 1443:30 FSM.scala 1445:27]
  wire [11:0] _GEN_1671 = _T_227 ? _L1_rd_addr_7_T_1 : _GEN_1660; // @[FSM.scala 1443:30 FSM.scala 1445:27]
  wire [11:0] _GEN_1672 = _T_227 ? _L1_rd_addr_8_T_1 : _GEN_1661; // @[FSM.scala 1443:30 FSM.scala 1445:27]
  wire [11:0] _GEN_1673 = _T_227 ? _L1_rd_addr_9_T_1 : _GEN_1662; // @[FSM.scala 1443:30 FSM.scala 1445:27]
  wire [11:0] _GEN_1674 = _T_227 ? _L1_rd_addr_10_T_1 : _GEN_1663; // @[FSM.scala 1443:30 FSM.scala 1445:27]
  wire [11:0] _GEN_1675 = _T_227 ? _L1_rd_addr_11_T_1 : _GEN_1664; // @[FSM.scala 1443:30 FSM.scala 1445:27]
  wire [11:0] _GEN_1676 = _T_228 ? _L1_rd_addr_2_T_1 : _GEN_1666; // @[FSM.scala 1448:30 FSM.scala 1450:27]
  wire [11:0] _GEN_1677 = _T_228 ? _L1_rd_addr_3_T_1 : _GEN_1667; // @[FSM.scala 1448:30 FSM.scala 1450:27]
  wire [11:0] _GEN_1678 = _T_228 ? _L1_rd_addr_4_T_1 : _GEN_1668; // @[FSM.scala 1448:30 FSM.scala 1450:27]
  wire [11:0] _GEN_1679 = _T_228 ? _L1_rd_addr_5_T_1 : _GEN_1669; // @[FSM.scala 1448:30 FSM.scala 1450:27]
  wire [11:0] _GEN_1680 = _T_228 ? _L1_rd_addr_6_T_1 : _GEN_1670; // @[FSM.scala 1448:30 FSM.scala 1450:27]
  wire [11:0] _GEN_1681 = _T_228 ? _L1_rd_addr_7_T_1 : _GEN_1671; // @[FSM.scala 1448:30 FSM.scala 1450:27]
  wire [11:0] _GEN_1682 = _T_228 ? _L1_rd_addr_8_T_1 : _GEN_1672; // @[FSM.scala 1448:30 FSM.scala 1450:27]
  wire [11:0] _GEN_1683 = _T_228 ? _L1_rd_addr_9_T_1 : _GEN_1673; // @[FSM.scala 1448:30 FSM.scala 1450:27]
  wire [11:0] _GEN_1684 = _T_228 ? _L1_rd_addr_10_T_1 : _GEN_1674; // @[FSM.scala 1448:30 FSM.scala 1450:27]
  wire [11:0] _GEN_1685 = _T_228 ? _L1_rd_addr_11_T_1 : _GEN_1675; // @[FSM.scala 1448:30 FSM.scala 1450:27]
  wire [11:0] _GEN_1686 = _T_229 ? _L1_rd_addr_3_T_1 : _GEN_1677; // @[FSM.scala 1453:30 FSM.scala 1455:27]
  wire [11:0] _GEN_1687 = _T_229 ? _L1_rd_addr_4_T_1 : _GEN_1678; // @[FSM.scala 1453:30 FSM.scala 1455:27]
  wire [11:0] _GEN_1688 = _T_229 ? _L1_rd_addr_5_T_1 : _GEN_1679; // @[FSM.scala 1453:30 FSM.scala 1455:27]
  wire [11:0] _GEN_1689 = _T_229 ? _L1_rd_addr_6_T_1 : _GEN_1680; // @[FSM.scala 1453:30 FSM.scala 1455:27]
  wire [11:0] _GEN_1690 = _T_229 ? _L1_rd_addr_7_T_1 : _GEN_1681; // @[FSM.scala 1453:30 FSM.scala 1455:27]
  wire [11:0] _GEN_1691 = _T_229 ? _L1_rd_addr_8_T_1 : _GEN_1682; // @[FSM.scala 1453:30 FSM.scala 1455:27]
  wire [11:0] _GEN_1692 = _T_229 ? _L1_rd_addr_9_T_1 : _GEN_1683; // @[FSM.scala 1453:30 FSM.scala 1455:27]
  wire [11:0] _GEN_1693 = _T_229 ? _L1_rd_addr_10_T_1 : _GEN_1684; // @[FSM.scala 1453:30 FSM.scala 1455:27]
  wire [11:0] _GEN_1694 = _T_229 ? _L1_rd_addr_11_T_1 : _GEN_1685; // @[FSM.scala 1453:30 FSM.scala 1455:27]
  wire [11:0] _GEN_1695 = _T_230 ? _L1_rd_addr_4_T_1 : _GEN_1687; // @[FSM.scala 1458:30 FSM.scala 1460:27]
  wire [11:0] _GEN_1696 = _T_230 ? _L1_rd_addr_5_T_1 : _GEN_1688; // @[FSM.scala 1458:30 FSM.scala 1460:27]
  wire [11:0] _GEN_1697 = _T_230 ? _L1_rd_addr_6_T_1 : _GEN_1689; // @[FSM.scala 1458:30 FSM.scala 1460:27]
  wire [11:0] _GEN_1698 = _T_230 ? _L1_rd_addr_7_T_1 : _GEN_1690; // @[FSM.scala 1458:30 FSM.scala 1460:27]
  wire [11:0] _GEN_1699 = _T_230 ? _L1_rd_addr_8_T_1 : _GEN_1691; // @[FSM.scala 1458:30 FSM.scala 1460:27]
  wire [11:0] _GEN_1700 = _T_230 ? _L1_rd_addr_9_T_1 : _GEN_1692; // @[FSM.scala 1458:30 FSM.scala 1460:27]
  wire [11:0] _GEN_1701 = _T_230 ? _L1_rd_addr_10_T_1 : _GEN_1693; // @[FSM.scala 1458:30 FSM.scala 1460:27]
  wire [11:0] _GEN_1702 = _T_230 ? _L1_rd_addr_11_T_1 : _GEN_1694; // @[FSM.scala 1458:30 FSM.scala 1460:27]
  wire [11:0] _GEN_1703 = _T_231 ? _L1_rd_addr_5_T_1 : _GEN_1696; // @[FSM.scala 1463:30 FSM.scala 1465:27]
  wire [11:0] _GEN_1704 = _T_231 ? _L1_rd_addr_6_T_1 : _GEN_1697; // @[FSM.scala 1463:30 FSM.scala 1465:27]
  wire [11:0] _GEN_1705 = _T_231 ? _L1_rd_addr_7_T_1 : _GEN_1698; // @[FSM.scala 1463:30 FSM.scala 1465:27]
  wire [11:0] _GEN_1706 = _T_231 ? _L1_rd_addr_8_T_1 : _GEN_1699; // @[FSM.scala 1463:30 FSM.scala 1465:27]
  wire [11:0] _GEN_1707 = _T_231 ? _L1_rd_addr_9_T_1 : _GEN_1700; // @[FSM.scala 1463:30 FSM.scala 1465:27]
  wire [11:0] _GEN_1708 = _T_231 ? _L1_rd_addr_10_T_1 : _GEN_1701; // @[FSM.scala 1463:30 FSM.scala 1465:27]
  wire [11:0] _GEN_1709 = _T_231 ? _L1_rd_addr_11_T_1 : _GEN_1702; // @[FSM.scala 1463:30 FSM.scala 1465:27]
  wire [11:0] _GEN_1710 = _T_232 ? _L1_rd_addr_6_T_1 : _GEN_1704; // @[FSM.scala 1468:30 FSM.scala 1470:27]
  wire [11:0] _GEN_1711 = _T_232 ? _L1_rd_addr_7_T_1 : _GEN_1705; // @[FSM.scala 1468:30 FSM.scala 1470:27]
  wire [11:0] _GEN_1712 = _T_232 ? _L1_rd_addr_8_T_1 : _GEN_1706; // @[FSM.scala 1468:30 FSM.scala 1470:27]
  wire [11:0] _GEN_1713 = _T_232 ? _L1_rd_addr_9_T_1 : _GEN_1707; // @[FSM.scala 1468:30 FSM.scala 1470:27]
  wire [11:0] _GEN_1714 = _T_232 ? _L1_rd_addr_10_T_1 : _GEN_1708; // @[FSM.scala 1468:30 FSM.scala 1470:27]
  wire [11:0] _GEN_1715 = _T_232 ? _L1_rd_addr_11_T_1 : _GEN_1709; // @[FSM.scala 1468:30 FSM.scala 1470:27]
  wire [11:0] _GEN_1716 = _T_233 ? _L1_rd_addr_7_T_1 : _GEN_1711; // @[FSM.scala 1473:30 FSM.scala 1475:27]
  wire [11:0] _GEN_1717 = _T_233 ? _L1_rd_addr_8_T_1 : _GEN_1712; // @[FSM.scala 1473:30 FSM.scala 1475:27]
  wire [11:0] _GEN_1718 = _T_233 ? _L1_rd_addr_9_T_1 : _GEN_1713; // @[FSM.scala 1473:30 FSM.scala 1475:27]
  wire [11:0] _GEN_1719 = _T_233 ? _L1_rd_addr_10_T_1 : _GEN_1714; // @[FSM.scala 1473:30 FSM.scala 1475:27]
  wire [11:0] _GEN_1720 = _T_233 ? _L1_rd_addr_11_T_1 : _GEN_1715; // @[FSM.scala 1473:30 FSM.scala 1475:27]
  wire [11:0] _GEN_1721 = _T_234 ? _L1_rd_addr_8_T_1 : _GEN_1717; // @[FSM.scala 1478:30 FSM.scala 1480:27]
  wire [11:0] _GEN_1722 = _T_234 ? _L1_rd_addr_9_T_1 : _GEN_1718; // @[FSM.scala 1478:30 FSM.scala 1480:27]
  wire [11:0] _GEN_1723 = _T_234 ? _L1_rd_addr_10_T_1 : _GEN_1719; // @[FSM.scala 1478:30 FSM.scala 1480:27]
  wire [11:0] _GEN_1724 = _T_234 ? _L1_rd_addr_11_T_1 : _GEN_1720; // @[FSM.scala 1478:30 FSM.scala 1480:27]
  wire [11:0] _GEN_1725 = _T_235 ? _L1_rd_addr_9_T_1 : _GEN_1722; // @[FSM.scala 1483:30 FSM.scala 1485:27]
  wire [11:0] _GEN_1726 = _T_235 ? _L1_rd_addr_10_T_1 : _GEN_1723; // @[FSM.scala 1483:30 FSM.scala 1485:27]
  wire [11:0] _GEN_1727 = _T_235 ? _L1_rd_addr_11_T_1 : _GEN_1724; // @[FSM.scala 1483:30 FSM.scala 1485:27]
  wire [11:0] _GEN_1728 = _T_236 ? _L1_rd_addr_10_T_1 : _GEN_1726; // @[FSM.scala 1488:30 FSM.scala 1490:27]
  wire [11:0] _GEN_1729 = _T_236 ? _L1_rd_addr_11_T_1 : _GEN_1727; // @[FSM.scala 1488:30 FSM.scala 1490:27]
  wire [11:0] _GEN_1730 = _T_65 ? _L1_rd_addr_11_T_1 : _GEN_1729; // @[FSM.scala 1493:30 FSM.scala 1495:27]
  wire [5:0] _FC_temp_wrAddr_T_1 = FC_temp_wrAddr + 6'h1; // @[FSM.scala 1505:48]
  wire [5:0] _GEN_1731 = _T_127 ? 6'h0 : _FC_temp_wrAddr_T_1; // @[FSM.scala 1500:33 FSM.scala 1501:28 FSM.scala 1505:30]
  wire [5:0] _GEN_1733 = _T_240 ? _GEN_1731 : _GEN_1576; // @[FSM.scala 1499:50]
  wire  _GEN_1734 = _T_240 | FC_temp_wrEna; // @[FSM.scala 1499:50 FSM.scala 96:38]
  wire [9:0] _GEN_1735 = _T_69 ? 10'h0 : _GEN_1567; // @[FSM.scala 1510:30 FSM.scala 1511:17]
  wire  _GEN_1737 = _T_69 ? 1'h0 : _GEN_1734; // @[FSM.scala 1510:30 FSM.scala 1513:25]
  wire [1:0] _GEN_1738 = _T_69 ? 2'h2 : _GEN_1566; // @[FSM.scala 1510:30 FSM.scala 1514:20]
  wire [9:0] _GEN_1739 = fc_state == 2'h1 ? _GEN_1735 : _GEN_1556; // @[FSM.scala 1338:29]
  wire [6:0] _GEN_1740 = fc_state == 2'h1 ? _GEN_1482 : count1; // @[FSM.scala 1338:29 FSM.scala 162:23]
  wire [2:0] _GEN_1741 = fc_state == 2'h1 ? _GEN_1579 : _GEN_1557; // @[FSM.scala 1338:29]
  wire [9:0] _GEN_1742 = fc_state == 2'h1 ? _GEN_1580 : _GEN_1559; // @[FSM.scala 1338:29]
  wire [5:0] _GEN_1743 = fc_state == 2'h1 ? _GEN_1581 : _GEN_1560; // @[FSM.scala 1338:29]
  wire [11:0] _GEN_1744 = fc_state == 2'h1 ? _GEN_1586 : _GEN_1558; // @[FSM.scala 1338:29]
  wire [7:0] _GEN_1745 = fc_state == 2'h1 ? _GEN_729 : PEArray_ctrl_2_gru_out_width; // @[FSM.scala 1338:29 FSM.scala 64:28]
  wire [1:0] _GEN_1746 = fc_state == 2'h1 ? _GEN_1574 : _GEN_1561; // @[FSM.scala 1338:29]
  wire [3:0] _GEN_1747 = fc_state == 2'h1 ? _GEN_1575 : _GEN_1562; // @[FSM.scala 1338:29]
  wire [5:0] _GEN_1748 = fc_state == 2'h1 ? _GEN_1733 : FC_temp_wrAddr; // @[FSM.scala 1338:29 FSM.scala 97:38]
  wire [1:0] _GEN_1749 = fc_state == 2'h1 ? _GEN_1577 : BN_Unit_ctrl; // @[FSM.scala 1338:29 FSM.scala 69:28]
  wire [1:0] _GEN_1750 = fc_state == 2'h1 ? _GEN_1578 : Activation_ctrl; // @[FSM.scala 1338:29 FSM.scala 75:32]
  wire [11:0] _GEN_1751 = fc_state == 2'h1 ? _GEN_1584 : _GEN_1563; // @[FSM.scala 1338:29]
  wire [11:0] _GEN_1752 = fc_state == 2'h1 ? _GEN_1585 : _GEN_1564; // @[FSM.scala 1338:29]
  wire [11:0] _GEN_1753 = fc_state == 2'h1 ? _GEN_1653 : L1_rd_addr_0; // @[FSM.scala 1338:29 FSM.scala 60:28]
  wire [11:0] _GEN_1754 = fc_state == 2'h1 ? _GEN_1665 : L1_rd_addr_1; // @[FSM.scala 1338:29 FSM.scala 60:28]
  wire [11:0] _GEN_1755 = fc_state == 2'h1 ? _GEN_1676 : L1_rd_addr_2; // @[FSM.scala 1338:29 FSM.scala 60:28]
  wire [11:0] _GEN_1756 = fc_state == 2'h1 ? _GEN_1686 : L1_rd_addr_3; // @[FSM.scala 1338:29 FSM.scala 60:28]
  wire [11:0] _GEN_1757 = fc_state == 2'h1 ? _GEN_1695 : L1_rd_addr_4; // @[FSM.scala 1338:29 FSM.scala 60:28]
  wire [11:0] _GEN_1758 = fc_state == 2'h1 ? _GEN_1703 : L1_rd_addr_5; // @[FSM.scala 1338:29 FSM.scala 60:28]
  wire [11:0] _GEN_1759 = fc_state == 2'h1 ? _GEN_1710 : L1_rd_addr_6; // @[FSM.scala 1338:29 FSM.scala 60:28]
  wire [11:0] _GEN_1760 = fc_state == 2'h1 ? _GEN_1716 : L1_rd_addr_7; // @[FSM.scala 1338:29 FSM.scala 60:28]
  wire [11:0] _GEN_1761 = fc_state == 2'h1 ? _GEN_1721 : L1_rd_addr_8; // @[FSM.scala 1338:29 FSM.scala 60:28]
  wire [11:0] _GEN_1762 = fc_state == 2'h1 ? _GEN_1725 : L1_rd_addr_9; // @[FSM.scala 1338:29 FSM.scala 60:28]
  wire [11:0] _GEN_1763 = fc_state == 2'h1 ? _GEN_1728 : L1_rd_addr_10; // @[FSM.scala 1338:29 FSM.scala 60:28]
  wire [11:0] _GEN_1764 = fc_state == 2'h1 ? _GEN_1730 : L1_rd_addr_11; // @[FSM.scala 1338:29 FSM.scala 60:28]
  wire  _GEN_1765 = fc_state == 2'h1 ? _GEN_1737 : FC_temp_wrEna; // @[FSM.scala 1338:29 FSM.scala 96:38]
  wire [1:0] _GEN_1766 = fc_state == 2'h1 ? _GEN_1738 : _GEN_1566; // @[FSM.scala 1338:29]
  wire [9:0] _GEN_1767 = _T_257 ? _count_T_1 : _GEN_1739; // @[FSM.scala 1518:29 FSM.scala 1519:17]
  wire [2:0] _GEN_1768 = _T_3 ? 3'h3 : _GEN_1741; // @[FSM.scala 1522:28 FSM.scala 1524:35]
  wire [11:0] _GEN_1769 = _T_3 ? 12'hfff : _GEN_1744; // @[FSM.scala 1522:28 FSM.scala 1525:32]
  wire [9:0] _GEN_1770 = _T_3 ? 10'h7 : _GEN_1742; // @[FSM.scala 1522:28 FSM.scala 1526:33]
  wire [5:0] _GEN_1771 = _T_3 ? 6'hf : _GEN_1743; // @[FSM.scala 1522:28 FSM.scala 1527:35]
  wire [1:0] _GEN_1772 = _T_3 ? 2'h2 : _GEN_1746; // @[FSM.scala 1522:28 FSM.scala 1529:30]
  wire [3:0] _GEN_1773 = _T_3 ? 4'h0 : _GEN_1747; // @[FSM.scala 1522:28 FSM.scala 1530:26]
  wire [11:0] _GEN_1774 = _T_5 ? 12'h0 : _GEN_1751; // @[FSM.scala 1532:28 FSM.scala 1534:34]
  wire [11:0] _GEN_1775 = _T_5 ? 12'h0 : _GEN_1752; // @[FSM.scala 1532:28 FSM.scala 1534:34]
  wire [11:0] _GEN_1776 = _T_5 ? 12'h0 : _GEN_1769; // @[FSM.scala 1532:28 FSM.scala 1534:34]
  wire [2:0] _GEN_1777 = _T_48 ? 3'h0 : FC_temp_to_PE_control; // @[FSM.scala 1537:28 FSM.scala 1538:33 FSM.scala 94:38]
  wire [2:0] _FC_temp_to_PE_control_T_1 = FC_temp_to_PE_control + 3'h1; // @[FSM.scala 1542:58]
  wire [2:0] _GEN_1778 = _T_85 ? _FC_temp_to_PE_control_T_1 : _GEN_1777; // @[FSM.scala 1541:47 FSM.scala 1542:33]
  wire [9:0] _GEN_1779 = _T_56 ? 10'h0 : _GEN_1767; // @[FSM.scala 1544:29 FSM.scala 1545:17]
  wire [1:0] _GEN_1780 = _T_56 ? 2'h3 : _GEN_1766; // @[FSM.scala 1544:29 FSM.scala 1546:20]
  wire [9:0] _GEN_1781 = fc_state == 2'h2 ? _GEN_1779 : _GEN_1739; // @[FSM.scala 1517:29]
  wire [2:0] _GEN_1782 = fc_state == 2'h2 ? _GEN_1768 : _GEN_1741; // @[FSM.scala 1517:29]
  wire [11:0] _GEN_1783 = fc_state == 2'h2 ? _GEN_1776 : _GEN_1744; // @[FSM.scala 1517:29]
  wire [9:0] _GEN_1784 = fc_state == 2'h2 ? _GEN_1770 : _GEN_1742; // @[FSM.scala 1517:29]
  wire [5:0] _GEN_1785 = fc_state == 2'h2 ? _GEN_1771 : _GEN_1743; // @[FSM.scala 1517:29]
  wire [1:0] _GEN_1786 = fc_state == 2'h2 ? _GEN_1772 : _GEN_1746; // @[FSM.scala 1517:29]
  wire [3:0] _GEN_1787 = fc_state == 2'h2 ? _GEN_1773 : _GEN_1747; // @[FSM.scala 1517:29]
  wire [11:0] _GEN_1788 = fc_state == 2'h2 ? _GEN_1774 : _GEN_1751; // @[FSM.scala 1517:29]
  wire [11:0] _GEN_1789 = fc_state == 2'h2 ? _GEN_1775 : _GEN_1752; // @[FSM.scala 1517:29]
  wire [2:0] _GEN_1790 = fc_state == 2'h2 ? _GEN_1778 : FC_temp_to_PE_control; // @[FSM.scala 1517:29 FSM.scala 94:38]
  wire [1:0] _GEN_1791 = fc_state == 2'h2 ? _GEN_1780 : _GEN_1766; // @[FSM.scala 1517:29]
  wire [9:0] _GEN_1792 = _T_206 ? _count_T_1 : _GEN_1781; // @[FSM.scala 1551:30 FSM.scala 1552:17]
  wire [6:0] _GEN_1793 = count1 != 7'hb ? _count1_T_1 : 7'h0; // @[FSM.scala 1555:30 FSM.scala 1556:18 FSM.scala 1558:18]
  wire [2:0] _GEN_1794 = _T_3 ? 3'h4 : _GEN_1782; // @[FSM.scala 1561:28 FSM.scala 1563:35]
  wire [9:0] _GEN_1795 = _T_3 ? 10'h47 : _GEN_1784; // @[FSM.scala 1561:28 FSM.scala 1564:33]
  wire [5:0] _GEN_1796 = _T_3 ? 6'hf : _GEN_1785; // @[FSM.scala 1561:28 FSM.scala 1565:35]
  wire [11:0] _GEN_1797 = _T_3 ? 12'h800 : _GEN_1783; // @[FSM.scala 1561:28 FSM.scala 1566:32]
  wire [7:0] _GEN_1798 = _T_3 ? 8'hc : _GEN_1745; // @[FSM.scala 1561:28 FSM.scala 1567:41]
  wire [1:0] _GEN_1799 = _T_3 ? 2'h0 : _GEN_1786; // @[FSM.scala 1561:28 FSM.scala 1570:30]
  wire [3:0] _GEN_1800 = _T_3 ? 4'h0 : _GEN_1787; // @[FSM.scala 1561:28 FSM.scala 1571:26]
  wire [5:0] _GEN_1801 = _T_3 ? 6'h0 : _GEN_1748; // @[FSM.scala 1561:28 FSM.scala 1574:26]
  wire [1:0] _GEN_1802 = _T_3 ? 2'h0 : _GEN_1749; // @[FSM.scala 1561:28 FSM.scala 1575:24]
  wire [1:0] _GEN_1803 = _T_3 ? 2'h0 : _GEN_1750; // @[FSM.scala 1561:28 FSM.scala 1576:27]
  wire [2:0] _GEN_1804 = _T_39 ? 3'h4 : _GEN_1794; // @[FSM.scala 1580:48 FSM.scala 1581:35]
  wire [9:0] _GEN_1805 = _T_39 ? 10'h47 : _GEN_1795; // @[FSM.scala 1580:48 FSM.scala 1582:33]
  wire [5:0] _GEN_1806 = _T_39 ? 6'hf : _GEN_1796; // @[FSM.scala 1580:48 FSM.scala 1583:35]
  wire [11:0] _GEN_1807 = _T_39 ? {{1'd0}, PEArray_ctrl_2_mask[11:1]} : _GEN_1797; // @[FSM.scala 1580:48 FSM.scala 1584:32]
  wire [7:0] _GEN_1808 = _T_39 ? 8'hc : _GEN_1798; // @[FSM.scala 1580:48 FSM.scala 1585:41]
  wire [11:0] _GEN_1809 = _T_40 ? 12'h0 : _GEN_1788; // @[FSM.scala 1587:29 FSM.scala 1589:34]
  wire [11:0] _GEN_1810 = _T_40 ? 12'h0 : _GEN_1789; // @[FSM.scala 1587:29 FSM.scala 1589:34]
  wire [11:0] _GEN_1811 = _T_40 ? 12'h0 : _GEN_1807; // @[FSM.scala 1587:29 FSM.scala 1589:34]
  wire [11:0] _GEN_1812 = _T_5 ? _L1_rd_addr_0_T_1 : _GEN_1753; // @[FSM.scala 1594:28 FSM.scala 1596:27]
  wire [11:0] _GEN_1813 = _T_48 ? _L1_rd_addr_0_T_1 : _GEN_1812; // @[FSM.scala 1599:28 FSM.scala 1601:27]
  wire [11:0] _GEN_1814 = _T_48 ? _L1_rd_addr_1_T_1 : _GEN_1754; // @[FSM.scala 1599:28 FSM.scala 1601:27]
  wire [11:0] _GEN_1815 = _T_49 ? _L1_rd_addr_0_T_1 : _GEN_1813; // @[FSM.scala 1604:28 FSM.scala 1606:27]
  wire [11:0] _GEN_1816 = _T_49 ? _L1_rd_addr_1_T_1 : _GEN_1814; // @[FSM.scala 1604:28 FSM.scala 1606:27]
  wire [11:0] _GEN_1817 = _T_49 ? _L1_rd_addr_2_T_1 : _GEN_1755; // @[FSM.scala 1604:28 FSM.scala 1606:27]
  wire [11:0] _GEN_1818 = _T_21 ? _L1_rd_addr_0_T_1 : _GEN_1815; // @[FSM.scala 1609:28 FSM.scala 1611:27]
  wire [11:0] _GEN_1819 = _T_21 ? _L1_rd_addr_1_T_1 : _GEN_1816; // @[FSM.scala 1609:28 FSM.scala 1611:27]
  wire [11:0] _GEN_1820 = _T_21 ? _L1_rd_addr_2_T_1 : _GEN_1817; // @[FSM.scala 1609:28 FSM.scala 1611:27]
  wire [11:0] _GEN_1821 = _T_21 ? _L1_rd_addr_3_T_1 : _GEN_1756; // @[FSM.scala 1609:28 FSM.scala 1611:27]
  wire [11:0] _GEN_1822 = _T_51 ? _L1_rd_addr_0_T_1 : _GEN_1818; // @[FSM.scala 1614:28 FSM.scala 1616:27]
  wire [11:0] _GEN_1823 = _T_51 ? _L1_rd_addr_1_T_1 : _GEN_1819; // @[FSM.scala 1614:28 FSM.scala 1616:27]
  wire [11:0] _GEN_1824 = _T_51 ? _L1_rd_addr_2_T_1 : _GEN_1820; // @[FSM.scala 1614:28 FSM.scala 1616:27]
  wire [11:0] _GEN_1825 = _T_51 ? _L1_rd_addr_3_T_1 : _GEN_1821; // @[FSM.scala 1614:28 FSM.scala 1616:27]
  wire [11:0] _GEN_1826 = _T_51 ? _L1_rd_addr_4_T_1 : _GEN_1757; // @[FSM.scala 1614:28 FSM.scala 1616:27]
  wire [11:0] _GEN_1827 = _T_52 ? _L1_rd_addr_0_T_1 : _GEN_1822; // @[FSM.scala 1619:28 FSM.scala 1621:27]
  wire [11:0] _GEN_1828 = _T_52 ? _L1_rd_addr_1_T_1 : _GEN_1823; // @[FSM.scala 1619:28 FSM.scala 1621:27]
  wire [11:0] _GEN_1829 = _T_52 ? _L1_rd_addr_2_T_1 : _GEN_1824; // @[FSM.scala 1619:28 FSM.scala 1621:27]
  wire [11:0] _GEN_1830 = _T_52 ? _L1_rd_addr_3_T_1 : _GEN_1825; // @[FSM.scala 1619:28 FSM.scala 1621:27]
  wire [11:0] _GEN_1831 = _T_52 ? _L1_rd_addr_4_T_1 : _GEN_1826; // @[FSM.scala 1619:28 FSM.scala 1621:27]
  wire [11:0] _GEN_1832 = _T_52 ? _L1_rd_addr_5_T_1 : _GEN_1758; // @[FSM.scala 1619:28 FSM.scala 1621:27]
  wire [11:0] _GEN_1833 = _T_53 ? _L1_rd_addr_0_T_1 : _GEN_1827; // @[FSM.scala 1624:28 FSM.scala 1626:27]
  wire [11:0] _GEN_1834 = _T_53 ? _L1_rd_addr_1_T_1 : _GEN_1828; // @[FSM.scala 1624:28 FSM.scala 1626:27]
  wire [11:0] _GEN_1835 = _T_53 ? _L1_rd_addr_2_T_1 : _GEN_1829; // @[FSM.scala 1624:28 FSM.scala 1626:27]
  wire [11:0] _GEN_1836 = _T_53 ? _L1_rd_addr_3_T_1 : _GEN_1830; // @[FSM.scala 1624:28 FSM.scala 1626:27]
  wire [11:0] _GEN_1837 = _T_53 ? _L1_rd_addr_4_T_1 : _GEN_1831; // @[FSM.scala 1624:28 FSM.scala 1626:27]
  wire [11:0] _GEN_1838 = _T_53 ? _L1_rd_addr_5_T_1 : _GEN_1832; // @[FSM.scala 1624:28 FSM.scala 1626:27]
  wire [11:0] _GEN_1839 = _T_53 ? _L1_rd_addr_6_T_1 : _GEN_1759; // @[FSM.scala 1624:28 FSM.scala 1626:27]
  wire [11:0] _GEN_1840 = _T_54 ? _L1_rd_addr_0_T_1 : _GEN_1833; // @[FSM.scala 1629:28 FSM.scala 1631:27]
  wire [11:0] _GEN_1841 = _T_54 ? _L1_rd_addr_1_T_1 : _GEN_1834; // @[FSM.scala 1629:28 FSM.scala 1631:27]
  wire [11:0] _GEN_1842 = _T_54 ? _L1_rd_addr_2_T_1 : _GEN_1835; // @[FSM.scala 1629:28 FSM.scala 1631:27]
  wire [11:0] _GEN_1843 = _T_54 ? _L1_rd_addr_3_T_1 : _GEN_1836; // @[FSM.scala 1629:28 FSM.scala 1631:27]
  wire [11:0] _GEN_1844 = _T_54 ? _L1_rd_addr_4_T_1 : _GEN_1837; // @[FSM.scala 1629:28 FSM.scala 1631:27]
  wire [11:0] _GEN_1845 = _T_54 ? _L1_rd_addr_5_T_1 : _GEN_1838; // @[FSM.scala 1629:28 FSM.scala 1631:27]
  wire [11:0] _GEN_1846 = _T_54 ? _L1_rd_addr_6_T_1 : _GEN_1839; // @[FSM.scala 1629:28 FSM.scala 1631:27]
  wire [11:0] _GEN_1847 = _T_54 ? _L1_rd_addr_7_T_1 : _GEN_1760; // @[FSM.scala 1629:28 FSM.scala 1631:27]
  wire [11:0] _GEN_1848 = _T_55 ? _L1_rd_addr_0_T_1 : _GEN_1840; // @[FSM.scala 1634:28 FSM.scala 1636:27]
  wire [11:0] _GEN_1849 = _T_55 ? _L1_rd_addr_1_T_1 : _GEN_1841; // @[FSM.scala 1634:28 FSM.scala 1636:27]
  wire [11:0] _GEN_1850 = _T_55 ? _L1_rd_addr_2_T_1 : _GEN_1842; // @[FSM.scala 1634:28 FSM.scala 1636:27]
  wire [11:0] _GEN_1851 = _T_55 ? _L1_rd_addr_3_T_1 : _GEN_1843; // @[FSM.scala 1634:28 FSM.scala 1636:27]
  wire [11:0] _GEN_1852 = _T_55 ? _L1_rd_addr_4_T_1 : _GEN_1844; // @[FSM.scala 1634:28 FSM.scala 1636:27]
  wire [11:0] _GEN_1853 = _T_55 ? _L1_rd_addr_5_T_1 : _GEN_1845; // @[FSM.scala 1634:28 FSM.scala 1636:27]
  wire [11:0] _GEN_1854 = _T_55 ? _L1_rd_addr_6_T_1 : _GEN_1846; // @[FSM.scala 1634:28 FSM.scala 1636:27]
  wire [11:0] _GEN_1855 = _T_55 ? _L1_rd_addr_7_T_1 : _GEN_1847; // @[FSM.scala 1634:28 FSM.scala 1636:27]
  wire [11:0] _GEN_1856 = _T_55 ? _L1_rd_addr_8_T_1 : _GEN_1761; // @[FSM.scala 1634:28 FSM.scala 1636:27]
  wire [11:0] _GEN_1857 = _T_56 ? _L1_rd_addr_0_T_1 : _GEN_1848; // @[FSM.scala 1639:29 FSM.scala 1641:27]
  wire [11:0] _GEN_1858 = _T_56 ? _L1_rd_addr_1_T_1 : _GEN_1849; // @[FSM.scala 1639:29 FSM.scala 1641:27]
  wire [11:0] _GEN_1859 = _T_56 ? _L1_rd_addr_2_T_1 : _GEN_1850; // @[FSM.scala 1639:29 FSM.scala 1641:27]
  wire [11:0] _GEN_1860 = _T_56 ? _L1_rd_addr_3_T_1 : _GEN_1851; // @[FSM.scala 1639:29 FSM.scala 1641:27]
  wire [11:0] _GEN_1861 = _T_56 ? _L1_rd_addr_4_T_1 : _GEN_1852; // @[FSM.scala 1639:29 FSM.scala 1641:27]
  wire [11:0] _GEN_1862 = _T_56 ? _L1_rd_addr_5_T_1 : _GEN_1853; // @[FSM.scala 1639:29 FSM.scala 1641:27]
  wire [11:0] _GEN_1863 = _T_56 ? _L1_rd_addr_6_T_1 : _GEN_1854; // @[FSM.scala 1639:29 FSM.scala 1641:27]
  wire [11:0] _GEN_1864 = _T_56 ? _L1_rd_addr_7_T_1 : _GEN_1855; // @[FSM.scala 1639:29 FSM.scala 1641:27]
  wire [11:0] _GEN_1865 = _T_56 ? _L1_rd_addr_8_T_1 : _GEN_1856; // @[FSM.scala 1639:29 FSM.scala 1641:27]
  wire [11:0] _GEN_1866 = _T_56 ? _L1_rd_addr_9_T_1 : _GEN_1762; // @[FSM.scala 1639:29 FSM.scala 1641:27]
  wire [11:0] _GEN_1867 = _T_57 ? _L1_rd_addr_0_T_1 : _GEN_1857; // @[FSM.scala 1644:29 FSM.scala 1646:27]
  wire [11:0] _GEN_1868 = _T_57 ? _L1_rd_addr_1_T_1 : _GEN_1858; // @[FSM.scala 1644:29 FSM.scala 1646:27]
  wire [11:0] _GEN_1869 = _T_57 ? _L1_rd_addr_2_T_1 : _GEN_1859; // @[FSM.scala 1644:29 FSM.scala 1646:27]
  wire [11:0] _GEN_1870 = _T_57 ? _L1_rd_addr_3_T_1 : _GEN_1860; // @[FSM.scala 1644:29 FSM.scala 1646:27]
  wire [11:0] _GEN_1871 = _T_57 ? _L1_rd_addr_4_T_1 : _GEN_1861; // @[FSM.scala 1644:29 FSM.scala 1646:27]
  wire [11:0] _GEN_1872 = _T_57 ? _L1_rd_addr_5_T_1 : _GEN_1862; // @[FSM.scala 1644:29 FSM.scala 1646:27]
  wire [11:0] _GEN_1873 = _T_57 ? _L1_rd_addr_6_T_1 : _GEN_1863; // @[FSM.scala 1644:29 FSM.scala 1646:27]
  wire [11:0] _GEN_1874 = _T_57 ? _L1_rd_addr_7_T_1 : _GEN_1864; // @[FSM.scala 1644:29 FSM.scala 1646:27]
  wire [11:0] _GEN_1875 = _T_57 ? _L1_rd_addr_8_T_1 : _GEN_1865; // @[FSM.scala 1644:29 FSM.scala 1646:27]
  wire [11:0] _GEN_1876 = _T_57 ? _L1_rd_addr_9_T_1 : _GEN_1866; // @[FSM.scala 1644:29 FSM.scala 1646:27]
  wire [11:0] _GEN_1877 = _T_57 ? _L1_rd_addr_10_T_1 : _GEN_1763; // @[FSM.scala 1644:29 FSM.scala 1646:27]
  wire [11:0] _GEN_1878 = _T_110 & count <= 10'h47 ? _L1_rd_addr_0_T_1 : _GEN_1867; // @[FSM.scala 1649:49 FSM.scala 1651:27]
  wire [11:0] _GEN_1879 = _T_110 & count <= 10'h47 ? _L1_rd_addr_1_T_1 : _GEN_1868; // @[FSM.scala 1649:49 FSM.scala 1651:27]
  wire [11:0] _GEN_1880 = _T_110 & count <= 10'h47 ? _L1_rd_addr_2_T_1 : _GEN_1869; // @[FSM.scala 1649:49 FSM.scala 1651:27]
  wire [11:0] _GEN_1881 = _T_110 & count <= 10'h47 ? _L1_rd_addr_3_T_1 : _GEN_1870; // @[FSM.scala 1649:49 FSM.scala 1651:27]
  wire [11:0] _GEN_1882 = _T_110 & count <= 10'h47 ? _L1_rd_addr_4_T_1 : _GEN_1871; // @[FSM.scala 1649:49 FSM.scala 1651:27]
  wire [11:0] _GEN_1883 = _T_110 & count <= 10'h47 ? _L1_rd_addr_5_T_1 : _GEN_1872; // @[FSM.scala 1649:49 FSM.scala 1651:27]
  wire [11:0] _GEN_1884 = _T_110 & count <= 10'h47 ? _L1_rd_addr_6_T_1 : _GEN_1873; // @[FSM.scala 1649:49 FSM.scala 1651:27]
  wire [11:0] _GEN_1885 = _T_110 & count <= 10'h47 ? _L1_rd_addr_7_T_1 : _GEN_1874; // @[FSM.scala 1649:49 FSM.scala 1651:27]
  wire [11:0] _GEN_1886 = _T_110 & count <= 10'h47 ? _L1_rd_addr_8_T_1 : _GEN_1875; // @[FSM.scala 1649:49 FSM.scala 1651:27]
  wire [11:0] _GEN_1887 = _T_110 & count <= 10'h47 ? _L1_rd_addr_9_T_1 : _GEN_1876; // @[FSM.scala 1649:49 FSM.scala 1651:27]
  wire [11:0] _GEN_1888 = _T_110 & count <= 10'h47 ? _L1_rd_addr_10_T_1 : _GEN_1877; // @[FSM.scala 1649:49 FSM.scala 1651:27]
  wire [11:0] _GEN_1889 = _T_110 & count <= 10'h47 ? _L1_rd_addr_11_T_1 : _GEN_1764; // @[FSM.scala 1649:49 FSM.scala 1651:27]
  wire [11:0] _GEN_1890 = count == 10'h48 ? _L1_rd_addr_1_T_1 : _GEN_1879; // @[FSM.scala 1654:29 FSM.scala 1656:27]
  wire [11:0] _GEN_1891 = count == 10'h48 ? _L1_rd_addr_2_T_1 : _GEN_1880; // @[FSM.scala 1654:29 FSM.scala 1656:27]
  wire [11:0] _GEN_1892 = count == 10'h48 ? _L1_rd_addr_3_T_1 : _GEN_1881; // @[FSM.scala 1654:29 FSM.scala 1656:27]
  wire [11:0] _GEN_1893 = count == 10'h48 ? _L1_rd_addr_4_T_1 : _GEN_1882; // @[FSM.scala 1654:29 FSM.scala 1656:27]
  wire [11:0] _GEN_1894 = count == 10'h48 ? _L1_rd_addr_5_T_1 : _GEN_1883; // @[FSM.scala 1654:29 FSM.scala 1656:27]
  wire [11:0] _GEN_1895 = count == 10'h48 ? _L1_rd_addr_6_T_1 : _GEN_1884; // @[FSM.scala 1654:29 FSM.scala 1656:27]
  wire [11:0] _GEN_1896 = count == 10'h48 ? _L1_rd_addr_7_T_1 : _GEN_1885; // @[FSM.scala 1654:29 FSM.scala 1656:27]
  wire [11:0] _GEN_1897 = count == 10'h48 ? _L1_rd_addr_8_T_1 : _GEN_1886; // @[FSM.scala 1654:29 FSM.scala 1656:27]
  wire [11:0] _GEN_1898 = count == 10'h48 ? _L1_rd_addr_9_T_1 : _GEN_1887; // @[FSM.scala 1654:29 FSM.scala 1656:27]
  wire [11:0] _GEN_1899 = count == 10'h48 ? _L1_rd_addr_10_T_1 : _GEN_1888; // @[FSM.scala 1654:29 FSM.scala 1656:27]
  wire [11:0] _GEN_1900 = count == 10'h48 ? _L1_rd_addr_11_T_1 : _GEN_1889; // @[FSM.scala 1654:29 FSM.scala 1656:27]
  wire [11:0] _GEN_1901 = count == 10'h49 ? _L1_rd_addr_2_T_1 : _GEN_1891; // @[FSM.scala 1659:29 FSM.scala 1661:27]
  wire [11:0] _GEN_1902 = count == 10'h49 ? _L1_rd_addr_3_T_1 : _GEN_1892; // @[FSM.scala 1659:29 FSM.scala 1661:27]
  wire [11:0] _GEN_1903 = count == 10'h49 ? _L1_rd_addr_4_T_1 : _GEN_1893; // @[FSM.scala 1659:29 FSM.scala 1661:27]
  wire [11:0] _GEN_1904 = count == 10'h49 ? _L1_rd_addr_5_T_1 : _GEN_1894; // @[FSM.scala 1659:29 FSM.scala 1661:27]
  wire [11:0] _GEN_1905 = count == 10'h49 ? _L1_rd_addr_6_T_1 : _GEN_1895; // @[FSM.scala 1659:29 FSM.scala 1661:27]
  wire [11:0] _GEN_1906 = count == 10'h49 ? _L1_rd_addr_7_T_1 : _GEN_1896; // @[FSM.scala 1659:29 FSM.scala 1661:27]
  wire [11:0] _GEN_1907 = count == 10'h49 ? _L1_rd_addr_8_T_1 : _GEN_1897; // @[FSM.scala 1659:29 FSM.scala 1661:27]
  wire [11:0] _GEN_1908 = count == 10'h49 ? _L1_rd_addr_9_T_1 : _GEN_1898; // @[FSM.scala 1659:29 FSM.scala 1661:27]
  wire [11:0] _GEN_1909 = count == 10'h49 ? _L1_rd_addr_10_T_1 : _GEN_1899; // @[FSM.scala 1659:29 FSM.scala 1661:27]
  wire [11:0] _GEN_1910 = count == 10'h49 ? _L1_rd_addr_11_T_1 : _GEN_1900; // @[FSM.scala 1659:29 FSM.scala 1661:27]
  wire [11:0] _GEN_1911 = count == 10'h4a ? _L1_rd_addr_3_T_1 : _GEN_1902; // @[FSM.scala 1664:29 FSM.scala 1666:27]
  wire [11:0] _GEN_1912 = count == 10'h4a ? _L1_rd_addr_4_T_1 : _GEN_1903; // @[FSM.scala 1664:29 FSM.scala 1666:27]
  wire [11:0] _GEN_1913 = count == 10'h4a ? _L1_rd_addr_5_T_1 : _GEN_1904; // @[FSM.scala 1664:29 FSM.scala 1666:27]
  wire [11:0] _GEN_1914 = count == 10'h4a ? _L1_rd_addr_6_T_1 : _GEN_1905; // @[FSM.scala 1664:29 FSM.scala 1666:27]
  wire [11:0] _GEN_1915 = count == 10'h4a ? _L1_rd_addr_7_T_1 : _GEN_1906; // @[FSM.scala 1664:29 FSM.scala 1666:27]
  wire [11:0] _GEN_1916 = count == 10'h4a ? _L1_rd_addr_8_T_1 : _GEN_1907; // @[FSM.scala 1664:29 FSM.scala 1666:27]
  wire [11:0] _GEN_1917 = count == 10'h4a ? _L1_rd_addr_9_T_1 : _GEN_1908; // @[FSM.scala 1664:29 FSM.scala 1666:27]
  wire [11:0] _GEN_1918 = count == 10'h4a ? _L1_rd_addr_10_T_1 : _GEN_1909; // @[FSM.scala 1664:29 FSM.scala 1666:27]
  wire [11:0] _GEN_1919 = count == 10'h4a ? _L1_rd_addr_11_T_1 : _GEN_1910; // @[FSM.scala 1664:29 FSM.scala 1666:27]
  wire [11:0] _GEN_1920 = count == 10'h4b ? _L1_rd_addr_4_T_1 : _GEN_1912; // @[FSM.scala 1669:29 FSM.scala 1671:27]
  wire [11:0] _GEN_1921 = count == 10'h4b ? _L1_rd_addr_5_T_1 : _GEN_1913; // @[FSM.scala 1669:29 FSM.scala 1671:27]
  wire [11:0] _GEN_1922 = count == 10'h4b ? _L1_rd_addr_6_T_1 : _GEN_1914; // @[FSM.scala 1669:29 FSM.scala 1671:27]
  wire [11:0] _GEN_1923 = count == 10'h4b ? _L1_rd_addr_7_T_1 : _GEN_1915; // @[FSM.scala 1669:29 FSM.scala 1671:27]
  wire [11:0] _GEN_1924 = count == 10'h4b ? _L1_rd_addr_8_T_1 : _GEN_1916; // @[FSM.scala 1669:29 FSM.scala 1671:27]
  wire [11:0] _GEN_1925 = count == 10'h4b ? _L1_rd_addr_9_T_1 : _GEN_1917; // @[FSM.scala 1669:29 FSM.scala 1671:27]
  wire [11:0] _GEN_1926 = count == 10'h4b ? _L1_rd_addr_10_T_1 : _GEN_1918; // @[FSM.scala 1669:29 FSM.scala 1671:27]
  wire [11:0] _GEN_1927 = count == 10'h4b ? _L1_rd_addr_11_T_1 : _GEN_1919; // @[FSM.scala 1669:29 FSM.scala 1671:27]
  wire [11:0] _GEN_1928 = count == 10'h4c ? _L1_rd_addr_5_T_1 : _GEN_1921; // @[FSM.scala 1674:29 FSM.scala 1676:27]
  wire [11:0] _GEN_1929 = count == 10'h4c ? _L1_rd_addr_6_T_1 : _GEN_1922; // @[FSM.scala 1674:29 FSM.scala 1676:27]
  wire [11:0] _GEN_1930 = count == 10'h4c ? _L1_rd_addr_7_T_1 : _GEN_1923; // @[FSM.scala 1674:29 FSM.scala 1676:27]
  wire [11:0] _GEN_1931 = count == 10'h4c ? _L1_rd_addr_8_T_1 : _GEN_1924; // @[FSM.scala 1674:29 FSM.scala 1676:27]
  wire [11:0] _GEN_1932 = count == 10'h4c ? _L1_rd_addr_9_T_1 : _GEN_1925; // @[FSM.scala 1674:29 FSM.scala 1676:27]
  wire [11:0] _GEN_1933 = count == 10'h4c ? _L1_rd_addr_10_T_1 : _GEN_1926; // @[FSM.scala 1674:29 FSM.scala 1676:27]
  wire [11:0] _GEN_1934 = count == 10'h4c ? _L1_rd_addr_11_T_1 : _GEN_1927; // @[FSM.scala 1674:29 FSM.scala 1676:27]
  wire [11:0] _GEN_1935 = count == 10'h4d ? _L1_rd_addr_6_T_1 : _GEN_1929; // @[FSM.scala 1679:29 FSM.scala 1681:27]
  wire [11:0] _GEN_1936 = count == 10'h4d ? _L1_rd_addr_7_T_1 : _GEN_1930; // @[FSM.scala 1679:29 FSM.scala 1681:27]
  wire [11:0] _GEN_1937 = count == 10'h4d ? _L1_rd_addr_8_T_1 : _GEN_1931; // @[FSM.scala 1679:29 FSM.scala 1681:27]
  wire [11:0] _GEN_1938 = count == 10'h4d ? _L1_rd_addr_9_T_1 : _GEN_1932; // @[FSM.scala 1679:29 FSM.scala 1681:27]
  wire [11:0] _GEN_1939 = count == 10'h4d ? _L1_rd_addr_10_T_1 : _GEN_1933; // @[FSM.scala 1679:29 FSM.scala 1681:27]
  wire [11:0] _GEN_1940 = count == 10'h4d ? _L1_rd_addr_11_T_1 : _GEN_1934; // @[FSM.scala 1679:29 FSM.scala 1681:27]
  wire [11:0] _GEN_1941 = count == 10'h4e ? _L1_rd_addr_7_T_1 : _GEN_1936; // @[FSM.scala 1684:29 FSM.scala 1686:27]
  wire [11:0] _GEN_1942 = count == 10'h4e ? _L1_rd_addr_8_T_1 : _GEN_1937; // @[FSM.scala 1684:29 FSM.scala 1686:27]
  wire [11:0] _GEN_1943 = count == 10'h4e ? _L1_rd_addr_9_T_1 : _GEN_1938; // @[FSM.scala 1684:29 FSM.scala 1686:27]
  wire [11:0] _GEN_1944 = count == 10'h4e ? _L1_rd_addr_10_T_1 : _GEN_1939; // @[FSM.scala 1684:29 FSM.scala 1686:27]
  wire [11:0] _GEN_1945 = count == 10'h4e ? _L1_rd_addr_11_T_1 : _GEN_1940; // @[FSM.scala 1684:29 FSM.scala 1686:27]
  wire [11:0] _GEN_1946 = count == 10'h4f ? _L1_rd_addr_8_T_1 : _GEN_1942; // @[FSM.scala 1689:29 FSM.scala 1691:27]
  wire [11:0] _GEN_1947 = count == 10'h4f ? _L1_rd_addr_9_T_1 : _GEN_1943; // @[FSM.scala 1689:29 FSM.scala 1691:27]
  wire [11:0] _GEN_1948 = count == 10'h4f ? _L1_rd_addr_10_T_1 : _GEN_1944; // @[FSM.scala 1689:29 FSM.scala 1691:27]
  wire [11:0] _GEN_1949 = count == 10'h4f ? _L1_rd_addr_11_T_1 : _GEN_1945; // @[FSM.scala 1689:29 FSM.scala 1691:27]
  wire [11:0] _GEN_1950 = count == 10'h50 ? _L1_rd_addr_9_T_1 : _GEN_1947; // @[FSM.scala 1694:29 FSM.scala 1696:27]
  wire [11:0] _GEN_1951 = count == 10'h50 ? _L1_rd_addr_10_T_1 : _GEN_1948; // @[FSM.scala 1694:29 FSM.scala 1696:27]
  wire [11:0] _GEN_1952 = count == 10'h50 ? _L1_rd_addr_11_T_1 : _GEN_1949; // @[FSM.scala 1694:29 FSM.scala 1696:27]
  wire [11:0] _GEN_1953 = count == 10'h51 ? _L1_rd_addr_10_T_1 : _GEN_1951; // @[FSM.scala 1699:29 FSM.scala 1701:27]
  wire [11:0] _GEN_1954 = count == 10'h51 ? _L1_rd_addr_11_T_1 : _GEN_1952; // @[FSM.scala 1699:29 FSM.scala 1701:27]
  wire [11:0] _GEN_1955 = count == 10'h52 ? _L1_rd_addr_11_T_1 : _GEN_1954; // @[FSM.scala 1704:29 FSM.scala 1706:27]
  wire [3:0] _Result_wrAddr_T_1 = Result_wrAddr + 4'h1; // @[FSM.scala 1716:46]
  wire [3:0] _GEN_1956 = _T_25 ? 4'h0 : _Result_wrAddr_T_1; // @[FSM.scala 1711:32 FSM.scala 1712:27 FSM.scala 1716:29]
  wire [3:0] _GEN_1958 = _T_124 & count <= 10'h55 ? _GEN_1956 : Result_wrAddr; // @[FSM.scala 1710:49 FSM.scala 100:38]
  wire  _GEN_1959 = _T_124 & count <= 10'h55 | Result_wrEna; // @[FSM.scala 1710:49 FSM.scala 99:38]
  wire [9:0] _GEN_1960 = count == 10'h56 ? 10'h0 : _GEN_1792; // @[FSM.scala 1721:29 FSM.scala 1722:17]
  wire [6:0] _GEN_1961 = count == 10'h56 ? 7'h0 : _GEN_1793; // @[FSM.scala 1721:29 FSM.scala 1723:18]
  wire  _GEN_1962 = count == 10'h56 ? 1'h0 : _GEN_1959; // @[FSM.scala 1721:29 FSM.scala 1724:24]
  wire [1:0] _GEN_1963 = count == 10'h56 ? 2'h0 : _GEN_1791; // @[FSM.scala 1721:29 FSM.scala 1725:20]
  wire [2:0] _GEN_1964 = count == 10'h56 ? 3'h0 : state; // @[FSM.scala 1721:29 FSM.scala 1726:17 FSM.scala 159:22]
  wire [9:0] _GEN_1965 = fc_state == 2'h3 ? _GEN_1960 : _GEN_1781; // @[FSM.scala 1550:29]
  wire [6:0] _GEN_1966 = fc_state == 2'h3 ? _GEN_1961 : _GEN_1740; // @[FSM.scala 1550:29]
  wire [2:0] _GEN_1967 = fc_state == 2'h3 ? _GEN_1804 : _GEN_1782; // @[FSM.scala 1550:29]
  wire [9:0] _GEN_1968 = fc_state == 2'h3 ? _GEN_1805 : _GEN_1784; // @[FSM.scala 1550:29]
  wire [5:0] _GEN_1969 = fc_state == 2'h3 ? _GEN_1806 : _GEN_1785; // @[FSM.scala 1550:29]
  wire [11:0] _GEN_1970 = fc_state == 2'h3 ? _GEN_1811 : _GEN_1783; // @[FSM.scala 1550:29]
  wire [7:0] _GEN_1971 = fc_state == 2'h3 ? _GEN_1808 : _GEN_1745; // @[FSM.scala 1550:29]
  wire [1:0] _GEN_1972 = fc_state == 2'h3 ? _GEN_1799 : _GEN_1786; // @[FSM.scala 1550:29]
  wire [3:0] _GEN_1973 = fc_state == 2'h3 ? _GEN_1800 : _GEN_1787; // @[FSM.scala 1550:29]
  wire [5:0] _GEN_1974 = fc_state == 2'h3 ? _GEN_1801 : _GEN_1748; // @[FSM.scala 1550:29]
  wire [1:0] _GEN_1975 = fc_state == 2'h3 ? _GEN_1802 : _GEN_1749; // @[FSM.scala 1550:29]
  wire [1:0] _GEN_1976 = fc_state == 2'h3 ? _GEN_1803 : _GEN_1750; // @[FSM.scala 1550:29]
  wire [11:0] _GEN_1977 = fc_state == 2'h3 ? _GEN_1809 : _GEN_1788; // @[FSM.scala 1550:29]
  wire [11:0] _GEN_1978 = fc_state == 2'h3 ? _GEN_1810 : _GEN_1789; // @[FSM.scala 1550:29]
  wire [11:0] _GEN_1979 = fc_state == 2'h3 ? _GEN_1878 : _GEN_1753; // @[FSM.scala 1550:29]
  wire [11:0] _GEN_1980 = fc_state == 2'h3 ? _GEN_1890 : _GEN_1754; // @[FSM.scala 1550:29]
  wire [11:0] _GEN_1981 = fc_state == 2'h3 ? _GEN_1901 : _GEN_1755; // @[FSM.scala 1550:29]
  wire [11:0] _GEN_1982 = fc_state == 2'h3 ? _GEN_1911 : _GEN_1756; // @[FSM.scala 1550:29]
  wire [11:0] _GEN_1983 = fc_state == 2'h3 ? _GEN_1920 : _GEN_1757; // @[FSM.scala 1550:29]
  wire [11:0] _GEN_1984 = fc_state == 2'h3 ? _GEN_1928 : _GEN_1758; // @[FSM.scala 1550:29]
  wire [11:0] _GEN_1985 = fc_state == 2'h3 ? _GEN_1935 : _GEN_1759; // @[FSM.scala 1550:29]
  wire [11:0] _GEN_1986 = fc_state == 2'h3 ? _GEN_1941 : _GEN_1760; // @[FSM.scala 1550:29]
  wire [11:0] _GEN_1987 = fc_state == 2'h3 ? _GEN_1946 : _GEN_1761; // @[FSM.scala 1550:29]
  wire [11:0] _GEN_1988 = fc_state == 2'h3 ? _GEN_1950 : _GEN_1762; // @[FSM.scala 1550:29]
  wire [11:0] _GEN_1989 = fc_state == 2'h3 ? _GEN_1953 : _GEN_1763; // @[FSM.scala 1550:29]
  wire [11:0] _GEN_1990 = fc_state == 2'h3 ? _GEN_1955 : _GEN_1764; // @[FSM.scala 1550:29]
  wire [3:0] _GEN_1991 = fc_state == 2'h3 ? _GEN_1958 : Result_wrAddr; // @[FSM.scala 1550:29 FSM.scala 100:38]
  wire  _GEN_1992 = fc_state == 2'h3 ? _GEN_1962 : Result_wrEna; // @[FSM.scala 1550:29 FSM.scala 99:38]
  wire [1:0] _GEN_1993 = fc_state == 2'h3 ? _GEN_1963 : _GEN_1791; // @[FSM.scala 1550:29]
  wire [2:0] _GEN_1994 = fc_state == 2'h3 ? _GEN_1964 : state; // @[FSM.scala 1550:29 FSM.scala 159:22]
  wire [9:0] _GEN_1995 = _T_255 ? _GEN_1965 : count; // @[Conditional.scala 39:67 FSM.scala 161:22]
  wire [2:0] _GEN_1996 = _T_255 ? _GEN_1967 : PEArray_ctrl_2_control; // @[Conditional.scala 39:67 FSM.scala 64:28]
  wire [11:0] _GEN_1997 = _T_255 ? _GEN_1970 : PEArray_ctrl_2_mask; // @[Conditional.scala 39:67 FSM.scala 64:28]
  wire [9:0] _GEN_1998 = _T_255 ? _GEN_1968 : PEArray_ctrl_2_count; // @[Conditional.scala 39:67 FSM.scala 64:28]
  wire [5:0] _GEN_1999 = _T_255 ? _GEN_1969 : PEArray_ctrl_2_L0index; // @[Conditional.scala 39:67 FSM.scala 64:28]
  wire [1:0] _GEN_2000 = _T_255 ? _GEN_1972 : PE_above_data_ctrl; // @[Conditional.scala 39:67 FSM.scala 74:35]
  wire [3:0] _GEN_2001 = _T_255 ? _GEN_1973 : PE_rd_data_mux; // @[Conditional.scala 39:67 FSM.scala 61:32]
  wire [11:0] _GEN_2002 = _T_255 ? _GEN_1977 : PEArray_ctrl_0_mask; // @[Conditional.scala 39:67 FSM.scala 64:28]
  wire [11:0] _GEN_2003 = _T_255 ? _GEN_1978 : PEArray_ctrl_1_mask; // @[Conditional.scala 39:67 FSM.scala 64:28]
  wire [2:0] _GEN_2004 = _T_255 ? _GEN_1565 : Ht_to_PE_control; // @[Conditional.scala 39:67 FSM.scala 77:36]
  wire [1:0] _GEN_2005 = _T_255 ? _GEN_1993 : fc_state; // @[Conditional.scala 39:67 FSM.scala 166:25]
  wire [6:0] _GEN_2006 = _T_255 ? _GEN_1966 : count1; // @[Conditional.scala 39:67 FSM.scala 162:23]
  wire [7:0] _GEN_2007 = _T_255 ? _GEN_1971 : PEArray_ctrl_2_gru_out_width; // @[Conditional.scala 39:67 FSM.scala 64:28]
  wire [5:0] _GEN_2008 = _T_255 ? _GEN_1974 : FC_temp_wrAddr; // @[Conditional.scala 39:67 FSM.scala 97:38]
  wire [1:0] _GEN_2009 = _T_255 ? _GEN_1975 : BN_Unit_ctrl; // @[Conditional.scala 39:67 FSM.scala 69:28]
  wire [1:0] _GEN_2010 = _T_255 ? _GEN_1976 : Activation_ctrl; // @[Conditional.scala 39:67 FSM.scala 75:32]
  wire [11:0] _GEN_2011 = _T_255 ? _GEN_1979 : L1_rd_addr_0; // @[Conditional.scala 39:67 FSM.scala 60:28]
  wire [11:0] _GEN_2012 = _T_255 ? _GEN_1980 : L1_rd_addr_1; // @[Conditional.scala 39:67 FSM.scala 60:28]
  wire [11:0] _GEN_2013 = _T_255 ? _GEN_1981 : L1_rd_addr_2; // @[Conditional.scala 39:67 FSM.scala 60:28]
  wire [11:0] _GEN_2014 = _T_255 ? _GEN_1982 : L1_rd_addr_3; // @[Conditional.scala 39:67 FSM.scala 60:28]
  wire [11:0] _GEN_2015 = _T_255 ? _GEN_1983 : L1_rd_addr_4; // @[Conditional.scala 39:67 FSM.scala 60:28]
  wire [11:0] _GEN_2016 = _T_255 ? _GEN_1984 : L1_rd_addr_5; // @[Conditional.scala 39:67 FSM.scala 60:28]
  wire [11:0] _GEN_2017 = _T_255 ? _GEN_1985 : L1_rd_addr_6; // @[Conditional.scala 39:67 FSM.scala 60:28]
  wire [11:0] _GEN_2018 = _T_255 ? _GEN_1986 : L1_rd_addr_7; // @[Conditional.scala 39:67 FSM.scala 60:28]
  wire [11:0] _GEN_2019 = _T_255 ? _GEN_1987 : L1_rd_addr_8; // @[Conditional.scala 39:67 FSM.scala 60:28]
  wire [11:0] _GEN_2020 = _T_255 ? _GEN_1988 : L1_rd_addr_9; // @[Conditional.scala 39:67 FSM.scala 60:28]
  wire [11:0] _GEN_2021 = _T_255 ? _GEN_1989 : L1_rd_addr_10; // @[Conditional.scala 39:67 FSM.scala 60:28]
  wire [11:0] _GEN_2022 = _T_255 ? _GEN_1990 : L1_rd_addr_11; // @[Conditional.scala 39:67 FSM.scala 60:28]
  wire  _GEN_2023 = _T_255 ? _GEN_1765 : FC_temp_wrEna; // @[Conditional.scala 39:67 FSM.scala 96:38]
  wire [2:0] _GEN_2024 = _T_255 ? _GEN_1790 : FC_temp_to_PE_control; // @[Conditional.scala 39:67 FSM.scala 94:38]
  wire [3:0] _GEN_2025 = _T_255 ? _GEN_1991 : Result_wrAddr; // @[Conditional.scala 39:67 FSM.scala 100:38]
  wire  _GEN_2026 = _T_255 ? _GEN_1992 : Result_wrEna; // @[Conditional.scala 39:67 FSM.scala 99:38]
  wire [2:0] _GEN_2027 = _T_255 ? _GEN_1994 : state; // @[Conditional.scala 39:67 FSM.scala 159:22]
  wire [9:0] _GEN_2028 = _T_77 ? _GEN_1532 : _GEN_1995; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_2029 = _T_77 ? _GEN_1487 : _GEN_1996; // @[Conditional.scala 39:67]
  wire [11:0] _GEN_2030 = _T_77 ? _GEN_1490 : _GEN_1997; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_2031 = _T_77 ? _GEN_1488 : _GEN_1998; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_2032 = _T_77 ? _GEN_1489 : _GEN_1999; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2033 = _T_77 ? _GEN_1492 : _GEN_2000; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_2034 = _T_77 ? _GEN_1493 : _GEN_2001; // @[Conditional.scala 39:67]
  wire [11:0] _GEN_2035 = _T_77 ? _GEN_1497 : _GEN_2002; // @[Conditional.scala 39:67]
  wire [11:0] _GEN_2036 = _T_77 ? _GEN_1498 : _GEN_2003; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_2037 = _T_77 ? _GEN_687 : _GEN_2004; // @[Conditional.scala 39:67]
  wire [11:0] _GEN_2038 = _T_77 ? _GEN_1499 : _GEN_2011; // @[Conditional.scala 39:67]
  wire [11:0] _GEN_2039 = _T_77 ? _GEN_1500 : _GEN_2012; // @[Conditional.scala 39:67]
  wire [11:0] _GEN_2040 = _T_77 ? _GEN_1501 : _GEN_2013; // @[Conditional.scala 39:67]
  wire [11:0] _GEN_2041 = _T_77 ? _GEN_1502 : _GEN_2014; // @[Conditional.scala 39:67]
  wire [11:0] _GEN_2042 = _T_77 ? _GEN_1503 : _GEN_2015; // @[Conditional.scala 39:67]
  wire [11:0] _GEN_2043 = _T_77 ? _GEN_1504 : _GEN_2016; // @[Conditional.scala 39:67]
  wire [11:0] _GEN_2044 = _T_77 ? _GEN_1505 : _GEN_2017; // @[Conditional.scala 39:67]
  wire [11:0] _GEN_2045 = _T_77 ? _GEN_1506 : _GEN_2018; // @[Conditional.scala 39:67]
  wire [11:0] _GEN_2046 = _T_77 ? _GEN_1507 : _GEN_2019; // @[Conditional.scala 39:67]
  wire [11:0] _GEN_2047 = _T_77 ? _GEN_1508 : _GEN_2020; // @[Conditional.scala 39:67]
  wire [11:0] _GEN_2048 = _T_77 ? _GEN_1509 : _GEN_2021; // @[Conditional.scala 39:67]
  wire [11:0] _GEN_2049 = _T_77 ? _GEN_1510 : _GEN_2022; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_2050 = _T_77 ? _GEN_1539 : gru_state; // @[Conditional.scala 39:67 FSM.scala 160:26]
  wire [6:0] _GEN_2051 = _T_77 ? _GEN_1486 : _GEN_2006; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_2052 = _T_77 ? _GEN_1491 : _GEN_2007; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_2053 = _T_77 ? _GEN_906 : Zt_wrAddr; // @[Conditional.scala 39:67 FSM.scala 83:36]
  wire [1:0] _GEN_2054 = _T_77 ? _GEN_1495 : _GEN_2009; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2055 = _T_77 ? _GEN_1496 : _GEN_2010; // @[Conditional.scala 39:67]
  wire  _GEN_2056 = _T_77 ? _GEN_911 : Zt_wrEna; // @[Conditional.scala 39:67 FSM.scala 82:36]
  wire [5:0] _GEN_2057 = _T_77 ? _GEN_1094 : Rt_wrAddr; // @[Conditional.scala 39:67 FSM.scala 86:36]
  wire  _GEN_2058 = _T_77 ? _GEN_1111 : Rt_wrEna; // @[Conditional.scala 39:67 FSM.scala 85:36]
  wire [5:0] _GEN_2059 = _T_77 ? _GEN_1294 : WhXt_wrAddr; // @[Conditional.scala 39:67 FSM.scala 89:36]
  wire  _GEN_2060 = _T_77 ? _GEN_1311 : WhXt_wrEna; // @[Conditional.scala 39:67 FSM.scala 88:36]
  wire [5:0] _GEN_2061 = _T_77 ? _GEN_1494 : Uhht_1_wrAddr; // @[Conditional.scala 39:67 FSM.scala 92:36]
  wire  _GEN_2062 = _T_77 ? _GEN_1511 : Uhht_1_wrEna; // @[Conditional.scala 39:67 FSM.scala 91:36]
  wire [5:0] _GEN_2063 = _T_77 ? _GEN_1533 : Zt_rdAddr; // @[Conditional.scala 39:67 FSM.scala 81:36]
  wire [5:0] _GEN_2064 = _T_77 ? _GEN_1534 : Rt_rdAddr; // @[Conditional.scala 39:67 FSM.scala 84:36]
  wire [5:0] _GEN_2065 = _T_77 ? _GEN_1535 : WhXt_rdAddr; // @[Conditional.scala 39:67 FSM.scala 87:36]
  wire [5:0] _GEN_2066 = _T_77 ? _GEN_1536 : Uhht_1_rdAddr; // @[Conditional.scala 39:67 FSM.scala 90:36]
  wire [5:0] _GEN_2067 = _T_77 ? _GEN_1537 : Ht_wrAddr; // @[Conditional.scala 39:67 FSM.scala 80:36]
  wire  _GEN_2068 = _T_77 ? _GEN_1538 : Ht_wrEna; // @[Conditional.scala 39:67 FSM.scala 79:36]
  wire [2:0] _GEN_2069 = _T_77 ? _GEN_1540 : _GEN_2027; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_2070 = _T_77 ? _GEN_1541 : gru_count; // @[Conditional.scala 39:67 FSM.scala 164:26]
  wire [1:0] _GEN_2071 = _T_77 ? fc_state : _GEN_2005; // @[Conditional.scala 39:67 FSM.scala 166:25]
  wire [5:0] _GEN_2072 = _T_77 ? FC_temp_wrAddr : _GEN_2008; // @[Conditional.scala 39:67 FSM.scala 97:38]
  wire  _GEN_2073 = _T_77 ? FC_temp_wrEna : _GEN_2023; // @[Conditional.scala 39:67 FSM.scala 96:38]
  wire [2:0] _GEN_2074 = _T_77 ? FC_temp_to_PE_control : _GEN_2024; // @[Conditional.scala 39:67 FSM.scala 94:38]
  wire [3:0] _GEN_2075 = _T_77 ? Result_wrAddr : _GEN_2025; // @[Conditional.scala 39:67 FSM.scala 100:38]
  wire  _GEN_2076 = _T_77 ? Result_wrEna : _GEN_2026; // @[Conditional.scala 39:67 FSM.scala 99:38]
  wire [9:0] _GEN_2077 = _T_32 ? _GEN_635 : _GEN_2028; // @[Conditional.scala 39:67]
  wire [6:0] _GEN_2078 = _T_32 ? _GEN_636 : _GEN_2051; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2093 = _T_32 ? _GEN_104 : _GEN_2033; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_2094 = _T_32 ? _GEN_334 : _GEN_2034; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_2133 = _T_32 ? _GEN_333 : read_index; // @[Conditional.scala 39:67 FSM.scala 165:27]
  wire [2:0] _GEN_2147 = _T_32 ? _GEN_638 : _GEN_2069; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_2150 = _T_32 ? Ht_to_PE_control : _GEN_2037; // @[Conditional.scala 39:67 FSM.scala 77:36]
  wire [3:0] _GEN_2151 = _T_32 ? gru_state : _GEN_2050; // @[Conditional.scala 39:67 FSM.scala 160:26]
  wire [5:0] _GEN_2153 = _T_32 ? Zt_wrAddr : _GEN_2053; // @[Conditional.scala 39:67 FSM.scala 83:36]
  wire [1:0] _GEN_2155 = _T_32 ? Activation_ctrl : _GEN_2055; // @[Conditional.scala 39:67 FSM.scala 75:32]
  wire  _GEN_2156 = _T_32 ? Zt_wrEna : _GEN_2056; // @[Conditional.scala 39:67 FSM.scala 82:36]
  wire [5:0] _GEN_2157 = _T_32 ? Rt_wrAddr : _GEN_2057; // @[Conditional.scala 39:67 FSM.scala 86:36]
  wire  _GEN_2158 = _T_32 ? Rt_wrEna : _GEN_2058; // @[Conditional.scala 39:67 FSM.scala 85:36]
  wire [5:0] _GEN_2159 = _T_32 ? WhXt_wrAddr : _GEN_2059; // @[Conditional.scala 39:67 FSM.scala 89:36]
  wire  _GEN_2160 = _T_32 ? WhXt_wrEna : _GEN_2060; // @[Conditional.scala 39:67 FSM.scala 88:36]
  wire [5:0] _GEN_2161 = _T_32 ? Uhht_1_wrAddr : _GEN_2061; // @[Conditional.scala 39:67 FSM.scala 92:36]
  wire  _GEN_2162 = _T_32 ? Uhht_1_wrEna : _GEN_2062; // @[Conditional.scala 39:67 FSM.scala 91:36]
  wire [5:0] _GEN_2163 = _T_32 ? Zt_rdAddr : _GEN_2063; // @[Conditional.scala 39:67 FSM.scala 81:36]
  wire [5:0] _GEN_2164 = _T_32 ? Rt_rdAddr : _GEN_2064; // @[Conditional.scala 39:67 FSM.scala 84:36]
  wire [5:0] _GEN_2165 = _T_32 ? WhXt_rdAddr : _GEN_2065; // @[Conditional.scala 39:67 FSM.scala 87:36]
  wire [5:0] _GEN_2166 = _T_32 ? Uhht_1_rdAddr : _GEN_2066; // @[Conditional.scala 39:67 FSM.scala 90:36]
  wire [5:0] _GEN_2167 = _T_32 ? Ht_wrAddr : _GEN_2067; // @[Conditional.scala 39:67 FSM.scala 80:36]
  wire  _GEN_2168 = _T_32 ? Ht_wrEna : _GEN_2068; // @[Conditional.scala 39:67 FSM.scala 79:36]
  wire [5:0] _GEN_2169 = _T_32 ? gru_count : _GEN_2070; // @[Conditional.scala 39:67 FSM.scala 164:26]
  wire [1:0] _GEN_2170 = _T_32 ? fc_state : _GEN_2071; // @[Conditional.scala 39:67 FSM.scala 166:25]
  wire [5:0] _GEN_2171 = _T_32 ? FC_temp_wrAddr : _GEN_2072; // @[Conditional.scala 39:67 FSM.scala 97:38]
  wire  _GEN_2172 = _T_32 ? FC_temp_wrEna : _GEN_2073; // @[Conditional.scala 39:67 FSM.scala 96:38]
  wire [2:0] _GEN_2173 = _T_32 ? FC_temp_to_PE_control : _GEN_2074; // @[Conditional.scala 39:67 FSM.scala 94:38]
  wire [3:0] _GEN_2174 = _T_32 ? Result_wrAddr : _GEN_2075; // @[Conditional.scala 39:67 FSM.scala 100:38]
  wire  _GEN_2175 = _T_32 ? Result_wrEna : _GEN_2076; // @[Conditional.scala 39:67 FSM.scala 99:38]
  wire  _GEN_2278 = _T_2 & _GEN_83; // @[Conditional.scala 39:67 FSM.scala 154:20]
  wire  _GEN_2279 = _T_2 ? _GEN_80 : Data_temp_used; // @[Conditional.scala 39:67 FSM.scala 105:31]
  wire  _GEN_2386 = _T ? Data_temp_used : _GEN_2279; // @[Conditional.scala 40:58 FSM.scala 105:31]
  assign io_Input_Ready = 1'h1; // @[FSM.scala 152:18]
  assign io_L1_wr_data = L1_wr_data; // @[FSM.scala 153:20]
  assign io_To_L1_control = _T ? 1'h0 : _GEN_2278; // @[Conditional.scala 40:58 FSM.scala 154:20]
  assign io_L1_rd_addr_0 = L1_rd_addr_0; // @[FSM.scala 110:21]
  assign io_L1_rd_addr_1 = L1_rd_addr_1; // @[FSM.scala 110:21]
  assign io_L1_rd_addr_2 = L1_rd_addr_2; // @[FSM.scala 110:21]
  assign io_L1_rd_addr_3 = L1_rd_addr_3; // @[FSM.scala 110:21]
  assign io_L1_rd_addr_4 = L1_rd_addr_4; // @[FSM.scala 110:21]
  assign io_L1_rd_addr_5 = L1_rd_addr_5; // @[FSM.scala 110:21]
  assign io_L1_rd_addr_6 = L1_rd_addr_6; // @[FSM.scala 110:21]
  assign io_L1_rd_addr_7 = L1_rd_addr_7; // @[FSM.scala 110:21]
  assign io_L1_rd_addr_8 = L1_rd_addr_8; // @[FSM.scala 110:21]
  assign io_L1_rd_addr_9 = L1_rd_addr_9; // @[FSM.scala 110:21]
  assign io_L1_rd_addr_10 = L1_rd_addr_10; // @[FSM.scala 110:21]
  assign io_L1_rd_addr_11 = L1_rd_addr_11; // @[FSM.scala 110:21]
  assign io_PE_rd_data_mux = PE_rd_data_mux; // @[FSM.scala 111:21]
  assign io_L1_wr_addr_0 = L1_wr_addr_0; // @[FSM.scala 112:21]
  assign io_L1_wr_addr_1 = L1_wr_addr_1; // @[FSM.scala 112:21]
  assign io_L1_wr_addr_2 = L1_wr_addr_2; // @[FSM.scala 112:21]
  assign io_L1_wr_addr_3 = L1_wr_addr_3; // @[FSM.scala 112:21]
  assign io_L1_wr_addr_4 = L1_wr_addr_4; // @[FSM.scala 112:21]
  assign io_L1_wr_addr_5 = L1_wr_addr_5; // @[FSM.scala 112:21]
  assign io_L1_wr_addr_6 = L1_wr_addr_6; // @[FSM.scala 112:21]
  assign io_L1_wr_addr_7 = L1_wr_addr_7; // @[FSM.scala 112:21]
  assign io_L1_wr_addr_8 = L1_wr_addr_8; // @[FSM.scala 112:21]
  assign io_L1_wr_addr_9 = L1_wr_addr_9; // @[FSM.scala 112:21]
  assign io_L1_wr_addr_10 = L1_wr_addr_10; // @[FSM.scala 112:21]
  assign io_L1_wr_addr_11 = L1_wr_addr_11; // @[FSM.scala 112:21]
  assign io_L1_wrEna_0 = L1_wrEna_0; // @[FSM.scala 113:21]
  assign io_L1_wrEna_1 = L1_wrEna_1; // @[FSM.scala 113:21]
  assign io_L1_wrEna_2 = L1_wrEna_2; // @[FSM.scala 113:21]
  assign io_L1_wrEna_3 = L1_wrEna_3; // @[FSM.scala 113:21]
  assign io_L1_wrEna_4 = L1_wrEna_4; // @[FSM.scala 113:21]
  assign io_L1_wrEna_5 = L1_wrEna_5; // @[FSM.scala 113:21]
  assign io_L1_wrEna_6 = L1_wrEna_6; // @[FSM.scala 113:21]
  assign io_L1_wrEna_7 = L1_wrEna_7; // @[FSM.scala 113:21]
  assign io_L1_wrEna_8 = L1_wrEna_8; // @[FSM.scala 113:21]
  assign io_L1_wrEna_9 = L1_wrEna_9; // @[FSM.scala 113:21]
  assign io_L1_wrEna_10 = L1_wrEna_10; // @[FSM.scala 113:21]
  assign io_L1_wrEna_11 = L1_wrEna_11; // @[FSM.scala 113:21]
  assign io_PEArray_ctrl_0_mask = PEArray_ctrl_0_mask; // @[FSM.scala 114:21]
  assign io_PEArray_ctrl_1_mask = PEArray_ctrl_1_mask; // @[FSM.scala 114:21]
  assign io_PEArray_ctrl_2_control = PEArray_ctrl_2_control; // @[FSM.scala 114:21]
  assign io_PEArray_ctrl_2_count = PEArray_ctrl_2_count; // @[FSM.scala 114:21]
  assign io_PEArray_ctrl_2_L0index = PEArray_ctrl_2_L0index; // @[FSM.scala 114:21]
  assign io_PEArray_ctrl_2_mask = PEArray_ctrl_2_mask; // @[FSM.scala 114:21]
  assign io_PEArray_ctrl_2_gru_out_width = PEArray_ctrl_2_gru_out_width; // @[FSM.scala 114:21]
  assign io_BNArray_ctrl_0 = BNArray_ctrl_0; // @[FSM.scala 115:21]
  assign io_BNArray_ctrl_1 = BNArray_ctrl_1; // @[FSM.scala 115:21]
  assign io_BNArray_ctrl_2 = BNArray_ctrl_2; // @[FSM.scala 115:21]
  assign io_BNArray_ctrl_3 = BNArray_ctrl_3; // @[FSM.scala 115:21]
  assign io_BNArray_ctrl_4 = BNArray_ctrl_4; // @[FSM.scala 115:21]
  assign io_BNArray_ctrl_5 = BNArray_ctrl_5; // @[FSM.scala 115:21]
  assign io_BNArray_ctrl_6 = BNArray_ctrl_6; // @[FSM.scala 115:21]
  assign io_BNArray_ctrl_7 = BNArray_ctrl_7; // @[FSM.scala 115:21]
  assign io_BNArray_ctrl_8 = BNArray_ctrl_8; // @[FSM.scala 115:21]
  assign io_BNArray_ctrl_9 = BNArray_ctrl_9; // @[FSM.scala 115:21]
  assign io_BNArray_ctrl_10 = BNArray_ctrl_10; // @[FSM.scala 115:21]
  assign io_BNArray_ctrl_11 = BNArray_ctrl_11; // @[FSM.scala 115:21]
  assign io_BN_Unit_ctrl = BN_Unit_ctrl; // @[FSM.scala 119:21]
  assign io_Relu6Array_ctrl_0 = Relu6Array_ctrl_0; // @[FSM.scala 123:21]
  assign io_Relu6Array_ctrl_1 = Relu6Array_ctrl_1; // @[FSM.scala 123:21]
  assign io_Relu6Array_ctrl_2 = Relu6Array_ctrl_2; // @[FSM.scala 123:21]
  assign io_Relu6Array_ctrl_3 = Relu6Array_ctrl_3; // @[FSM.scala 123:21]
  assign io_Relu6Array_ctrl_4 = Relu6Array_ctrl_4; // @[FSM.scala 123:21]
  assign io_Relu6Array_ctrl_5 = Relu6Array_ctrl_5; // @[FSM.scala 123:21]
  assign io_Relu6Array_ctrl_6 = Relu6Array_ctrl_6; // @[FSM.scala 123:21]
  assign io_Relu6Array_ctrl_7 = Relu6Array_ctrl_7; // @[FSM.scala 123:21]
  assign io_Relu6Array_ctrl_8 = Relu6Array_ctrl_8; // @[FSM.scala 123:21]
  assign io_Relu6Array_ctrl_9 = Relu6Array_ctrl_9; // @[FSM.scala 123:21]
  assign io_Relu6Array_ctrl_10 = Relu6Array_ctrl_10; // @[FSM.scala 123:21]
  assign io_Relu6Array_ctrl_11 = Relu6Array_ctrl_11; // @[FSM.scala 123:21]
  assign io_PE_above_data_ctrl = PE_above_data_ctrl; // @[FSM.scala 124:25]
  assign io_Activation_ctrl = Activation_ctrl; // @[FSM.scala 125:22]
  assign io_Ht_to_PE_control = Ht_to_PE_control; // @[FSM.scala 127:23]
  assign io_Ht_wrEna = Ht_wrEna; // @[FSM.scala 129:23]
  assign io_Ht_wrAddr = Ht_wrAddr; // @[FSM.scala 130:23]
  assign io_Zt_rdAddr = Zt_rdAddr; // @[FSM.scala 131:23]
  assign io_Zt_wrEna = Zt_wrEna; // @[FSM.scala 132:23]
  assign io_Zt_wrAddr = Zt_wrAddr; // @[FSM.scala 133:23]
  assign io_Rt_rdAddr = Rt_rdAddr; // @[FSM.scala 134:23]
  assign io_Rt_wrEna = Rt_wrEna; // @[FSM.scala 135:23]
  assign io_Rt_wrAddr = Rt_wrAddr; // @[FSM.scala 136:23]
  assign io_WhXt_rdAddr = WhXt_rdAddr; // @[FSM.scala 137:23]
  assign io_WhXt_wrEna = WhXt_wrEna; // @[FSM.scala 138:23]
  assign io_WhXt_wrAddr = WhXt_wrAddr; // @[FSM.scala 139:23]
  assign io_Uhht_1_rdAddr = Uhht_1_rdAddr; // @[FSM.scala 140:23]
  assign io_Uhht_1_wrEna = Uhht_1_wrEna; // @[FSM.scala 141:23]
  assign io_Uhht_1_wrAddr = Uhht_1_wrAddr; // @[FSM.scala 142:23]
  assign io_FC_temp_to_PE_control = FC_temp_to_PE_control; // @[FSM.scala 144:28]
  assign io_FC_temp_wrEna = FC_temp_wrEna; // @[FSM.scala 146:28]
  assign io_FC_temp_wrAddr = FC_temp_wrAddr; // @[FSM.scala 147:28]
  assign io_Result_wrEna = Result_wrEna; // @[FSM.scala 149:28]
  assign io_Result_wrAddr = Result_wrAddr; // @[FSM.scala 150:28]
  always @(posedge clock) begin
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          if (count >= 10'h1 & count <= 10'h31) begin // @[FSM.scala 241:46]
            L1_rd_addr_0 <= _L1_rd_addr_0_T_1; // @[FSM.scala 243:25]
          end else begin
            L1_rd_addr_0 <= _GEN_92;
          end
        end else if (_T_32) begin // @[Conditional.scala 39:67]
          L1_rd_addr_0 <= _GEN_321;
        end else begin
          L1_rd_addr_0 <= _GEN_2038;
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          if (count >= 10'h1 & count <= 10'h31) begin // @[FSM.scala 241:46]
            L1_rd_addr_1 <= _L1_rd_addr_1_T_1; // @[FSM.scala 243:25]
          end else begin
            L1_rd_addr_1 <= _GEN_93;
          end
        end else if (_T_32) begin // @[Conditional.scala 39:67]
          L1_rd_addr_1 <= _GEN_322;
        end else begin
          L1_rd_addr_1 <= _GEN_2039;
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          if (count >= 10'h1 & count <= 10'h31) begin // @[FSM.scala 241:46]
            L1_rd_addr_2 <= _L1_rd_addr_2_T_1; // @[FSM.scala 243:25]
          end else begin
            L1_rd_addr_2 <= _GEN_94;
          end
        end else if (_T_32) begin // @[Conditional.scala 39:67]
          L1_rd_addr_2 <= _GEN_323;
        end else begin
          L1_rd_addr_2 <= _GEN_2040;
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          if (count >= 10'h1 & count <= 10'h31) begin // @[FSM.scala 241:46]
            L1_rd_addr_3 <= _L1_rd_addr_3_T_1; // @[FSM.scala 243:25]
          end else begin
            L1_rd_addr_3 <= _GEN_95;
          end
        end else if (_T_32) begin // @[Conditional.scala 39:67]
          L1_rd_addr_3 <= _GEN_324;
        end else begin
          L1_rd_addr_3 <= _GEN_2041;
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          if (count >= 10'h1 & count <= 10'h31) begin // @[FSM.scala 241:46]
            L1_rd_addr_4 <= _L1_rd_addr_4_T_1; // @[FSM.scala 243:25]
          end else begin
            L1_rd_addr_4 <= _GEN_96;
          end
        end else if (_T_32) begin // @[Conditional.scala 39:67]
          L1_rd_addr_4 <= _GEN_325;
        end else begin
          L1_rd_addr_4 <= _GEN_2042;
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          if (count >= 10'h1 & count <= 10'h31) begin // @[FSM.scala 241:46]
            L1_rd_addr_5 <= _L1_rd_addr_5_T_1; // @[FSM.scala 243:25]
          end else begin
            L1_rd_addr_5 <= _GEN_97;
          end
        end else if (_T_32) begin // @[Conditional.scala 39:67]
          L1_rd_addr_5 <= _GEN_326;
        end else begin
          L1_rd_addr_5 <= _GEN_2043;
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          if (count >= 10'h1 & count <= 10'h31) begin // @[FSM.scala 241:46]
            L1_rd_addr_6 <= _L1_rd_addr_6_T_1; // @[FSM.scala 243:25]
          end else begin
            L1_rd_addr_6 <= _GEN_98;
          end
        end else if (_T_32) begin // @[Conditional.scala 39:67]
          L1_rd_addr_6 <= _GEN_327;
        end else begin
          L1_rd_addr_6 <= _GEN_2044;
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          if (count >= 10'h1 & count <= 10'h31) begin // @[FSM.scala 241:46]
            L1_rd_addr_7 <= _L1_rd_addr_7_T_1; // @[FSM.scala 243:25]
          end else begin
            L1_rd_addr_7 <= _GEN_99;
          end
        end else if (_T_32) begin // @[Conditional.scala 39:67]
          L1_rd_addr_7 <= _GEN_328;
        end else begin
          L1_rd_addr_7 <= _GEN_2045;
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          if (count >= 10'h1 & count <= 10'h31) begin // @[FSM.scala 241:46]
            L1_rd_addr_8 <= _L1_rd_addr_8_T_1; // @[FSM.scala 243:25]
          end else begin
            L1_rd_addr_8 <= _GEN_100;
          end
        end else if (_T_32) begin // @[Conditional.scala 39:67]
          L1_rd_addr_8 <= _GEN_329;
        end else begin
          L1_rd_addr_8 <= _GEN_2046;
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          if (count >= 10'h1 & count <= 10'h31) begin // @[FSM.scala 241:46]
            L1_rd_addr_9 <= _L1_rd_addr_9_T_1; // @[FSM.scala 243:25]
          end else begin
            L1_rd_addr_9 <= _GEN_101;
          end
        end else if (_T_32) begin // @[Conditional.scala 39:67]
          L1_rd_addr_9 <= _GEN_330;
        end else begin
          L1_rd_addr_9 <= _GEN_2047;
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          if (count >= 10'h1 & count <= 10'h31) begin // @[FSM.scala 241:46]
            L1_rd_addr_10 <= _L1_rd_addr_10_T_1; // @[FSM.scala 243:25]
          end else begin
            L1_rd_addr_10 <= _GEN_102;
          end
        end else if (_T_32) begin // @[Conditional.scala 39:67]
          L1_rd_addr_10 <= _GEN_331;
        end else begin
          L1_rd_addr_10 <= _GEN_2048;
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          if (count >= 10'h1 & count <= 10'h31) begin // @[FSM.scala 241:46]
            L1_rd_addr_11 <= _L1_rd_addr_11_T_1; // @[FSM.scala 243:25]
          end else begin
            L1_rd_addr_11 <= _GEN_103;
          end
        end else if (_T_32) begin // @[Conditional.scala 39:67]
          L1_rd_addr_11 <= _GEN_332;
        end else begin
          L1_rd_addr_11 <= _GEN_2049;
        end
      end
    end
    if (reset) begin // @[FSM.scala 61:32]
      PE_rd_data_mux <= 4'h0; // @[FSM.scala 61:32]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          PE_rd_data_mux <= _GEN_105;
        end else begin
          PE_rd_data_mux <= _GEN_2094;
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_2) begin // @[Conditional.scala 39:67]
        if (~Data_temp_used) begin // @[FSM.scala 179:39]
          if (count >= 10'h2 & count <= 10'hf) begin // @[FSM.scala 189:44]
            L1_wr_addr_0 <= _L1_wr_addr_0_T_1; // @[FSM.scala 192:27]
          end else begin
            L1_wr_addr_0 <= _GEN_4;
          end
        end
      end else if (_T_13) begin // @[Conditional.scala 39:67]
        if (count >= 10'h2c & count <= 10'h33) begin // @[FSM.scala 268:47]
          L1_wr_addr_0 <= _L1_wr_addr_0_T_1; // @[FSM.scala 270:23]
        end else begin
          L1_wr_addr_0 <= _GEN_194;
        end
      end else if (_T_32) begin // @[Conditional.scala 39:67]
        L1_wr_addr_0 <= _GEN_468;
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_2) begin // @[Conditional.scala 39:67]
        if (~Data_temp_used) begin // @[FSM.scala 179:39]
          if (count >= 10'h2 & count <= 10'hf) begin // @[FSM.scala 189:44]
            L1_wr_addr_1 <= _L1_wr_addr_1_T_1; // @[FSM.scala 192:27]
          end else begin
            L1_wr_addr_1 <= _GEN_6;
          end
        end
      end else if (_T_13) begin // @[Conditional.scala 39:67]
        if (count >= 10'h5 & count <= 10'h2b) begin // @[FSM.scala 256:46]
          L1_wr_addr_1 <= _GEN_171;
        end else begin
          L1_wr_addr_1 <= _GEN_126;
        end
      end else if (_T_32) begin // @[Conditional.scala 39:67]
        L1_wr_addr_1 <= _GEN_492;
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_2) begin // @[Conditional.scala 39:67]
        if (~Data_temp_used) begin // @[FSM.scala 179:39]
          if (count >= 10'h2 & count <= 10'hf) begin // @[FSM.scala 189:44]
            L1_wr_addr_2 <= _L1_wr_addr_2_T_1; // @[FSM.scala 192:27]
          end else begin
            L1_wr_addr_2 <= _GEN_8;
          end
        end
      end else if (_T_13) begin // @[Conditional.scala 39:67]
        if (count >= 10'h5 & count <= 10'h2b) begin // @[FSM.scala 256:46]
          L1_wr_addr_2 <= _GEN_172;
        end else begin
          L1_wr_addr_2 <= _GEN_130;
        end
      end else if (_T_32) begin // @[Conditional.scala 39:67]
        L1_wr_addr_2 <= _GEN_514;
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_2) begin // @[Conditional.scala 39:67]
        if (~Data_temp_used) begin // @[FSM.scala 179:39]
          if (count >= 10'h2 & count <= 10'hf) begin // @[FSM.scala 189:44]
            L1_wr_addr_3 <= _L1_wr_addr_3_T_1; // @[FSM.scala 192:27]
          end else begin
            L1_wr_addr_3 <= _GEN_10;
          end
        end
      end else if (_T_13) begin // @[Conditional.scala 39:67]
        if (count >= 10'h5 & count <= 10'h2b) begin // @[FSM.scala 256:46]
          L1_wr_addr_3 <= _GEN_173;
        end else begin
          L1_wr_addr_3 <= _GEN_134;
        end
      end else if (_T_32) begin // @[Conditional.scala 39:67]
        L1_wr_addr_3 <= _GEN_534;
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_2) begin // @[Conditional.scala 39:67]
        if (~Data_temp_used) begin // @[FSM.scala 179:39]
          if (count >= 10'h2 & count <= 10'hf) begin // @[FSM.scala 189:44]
            L1_wr_addr_4 <= _L1_wr_addr_4_T_1; // @[FSM.scala 192:27]
          end else begin
            L1_wr_addr_4 <= _GEN_12;
          end
        end
      end else if (_T_13) begin // @[Conditional.scala 39:67]
        if (count >= 10'h5 & count <= 10'h2b) begin // @[FSM.scala 256:46]
          L1_wr_addr_4 <= _GEN_174;
        end else begin
          L1_wr_addr_4 <= _GEN_138;
        end
      end else if (_T_32) begin // @[Conditional.scala 39:67]
        L1_wr_addr_4 <= _GEN_552;
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_2) begin // @[Conditional.scala 39:67]
        if (~Data_temp_used) begin // @[FSM.scala 179:39]
          if (count >= 10'h2 & count <= 10'hf) begin // @[FSM.scala 189:44]
            L1_wr_addr_5 <= _L1_wr_addr_5_T_1; // @[FSM.scala 192:27]
          end else begin
            L1_wr_addr_5 <= _GEN_14;
          end
        end
      end else if (_T_13) begin // @[Conditional.scala 39:67]
        if (count >= 10'h5 & count <= 10'h2b) begin // @[FSM.scala 256:46]
          L1_wr_addr_5 <= _GEN_175;
        end else begin
          L1_wr_addr_5 <= _GEN_142;
        end
      end else if (_T_32) begin // @[Conditional.scala 39:67]
        L1_wr_addr_5 <= _GEN_568;
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_2) begin // @[Conditional.scala 39:67]
        if (~Data_temp_used) begin // @[FSM.scala 179:39]
          if (count >= 10'h2 & count <= 10'hf) begin // @[FSM.scala 189:44]
            L1_wr_addr_6 <= _L1_wr_addr_6_T_1; // @[FSM.scala 192:27]
          end else begin
            L1_wr_addr_6 <= _GEN_16;
          end
        end
      end else if (_T_13) begin // @[Conditional.scala 39:67]
        if (count >= 10'h5 & count <= 10'h2b) begin // @[FSM.scala 256:46]
          L1_wr_addr_6 <= _GEN_176;
        end else begin
          L1_wr_addr_6 <= _GEN_146;
        end
      end else if (_T_32) begin // @[Conditional.scala 39:67]
        L1_wr_addr_6 <= _GEN_582;
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_2) begin // @[Conditional.scala 39:67]
        if (~Data_temp_used) begin // @[FSM.scala 179:39]
          if (count >= 10'h2 & count <= 10'hf) begin // @[FSM.scala 189:44]
            L1_wr_addr_7 <= _L1_wr_addr_7_T_1; // @[FSM.scala 192:27]
          end else begin
            L1_wr_addr_7 <= _GEN_18;
          end
        end
      end else if (_T_13) begin // @[Conditional.scala 39:67]
        if (count >= 10'h5 & count <= 10'h2b) begin // @[FSM.scala 256:46]
          L1_wr_addr_7 <= _GEN_177;
        end else begin
          L1_wr_addr_7 <= _GEN_150;
        end
      end else if (_T_32) begin // @[Conditional.scala 39:67]
        L1_wr_addr_7 <= _GEN_594;
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_2) begin // @[Conditional.scala 39:67]
        if (~Data_temp_used) begin // @[FSM.scala 179:39]
          if (count >= 10'h2 & count <= 10'hf) begin // @[FSM.scala 189:44]
            L1_wr_addr_8 <= _L1_wr_addr_8_T_1; // @[FSM.scala 192:27]
          end else begin
            L1_wr_addr_8 <= _GEN_20;
          end
        end
      end else if (_T_13) begin // @[Conditional.scala 39:67]
        if (count >= 10'h5 & count <= 10'h2b) begin // @[FSM.scala 256:46]
          L1_wr_addr_8 <= _GEN_178;
        end else begin
          L1_wr_addr_8 <= _GEN_154;
        end
      end else if (_T_32) begin // @[Conditional.scala 39:67]
        L1_wr_addr_8 <= _GEN_604;
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_2) begin // @[Conditional.scala 39:67]
        if (~Data_temp_used) begin // @[FSM.scala 179:39]
          if (count >= 10'h2 & count <= 10'hf) begin // @[FSM.scala 189:44]
            L1_wr_addr_9 <= _L1_wr_addr_9_T_1; // @[FSM.scala 192:27]
          end else begin
            L1_wr_addr_9 <= _GEN_22;
          end
        end
      end else if (_T_13) begin // @[Conditional.scala 39:67]
        if (count >= 10'h5 & count <= 10'h2b) begin // @[FSM.scala 256:46]
          L1_wr_addr_9 <= _GEN_179;
        end else begin
          L1_wr_addr_9 <= _GEN_158;
        end
      end else if (_T_32) begin // @[Conditional.scala 39:67]
        L1_wr_addr_9 <= _GEN_612;
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_2) begin // @[Conditional.scala 39:67]
        if (~Data_temp_used) begin // @[FSM.scala 179:39]
          if (count >= 10'h2 & count <= 10'hf) begin // @[FSM.scala 189:44]
            L1_wr_addr_10 <= _L1_wr_addr_10_T_1; // @[FSM.scala 192:27]
          end else begin
            L1_wr_addr_10 <= _GEN_24;
          end
        end
      end else if (_T_13) begin // @[Conditional.scala 39:67]
        if (count >= 10'h5 & count <= 10'h2b) begin // @[FSM.scala 256:46]
          L1_wr_addr_10 <= _GEN_180;
        end else begin
          L1_wr_addr_10 <= _GEN_162;
        end
      end else if (_T_32) begin // @[Conditional.scala 39:67]
        L1_wr_addr_10 <= _GEN_618;
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_2) begin // @[Conditional.scala 39:67]
        if (~Data_temp_used) begin // @[FSM.scala 179:39]
          if (count >= 10'h2 & count <= 10'hf) begin // @[FSM.scala 189:44]
            L1_wr_addr_11 <= _L1_wr_addr_11_T_1; // @[FSM.scala 192:27]
          end else begin
            L1_wr_addr_11 <= _GEN_26;
          end
        end
      end else if (_T_13) begin // @[Conditional.scala 39:67]
        if (count >= 10'h5 & count <= 10'h2b) begin // @[FSM.scala 256:46]
          L1_wr_addr_11 <= _GEN_181;
        end else begin
          L1_wr_addr_11 <= _GEN_166;
        end
      end else if (_T_32) begin // @[Conditional.scala 39:67]
        L1_wr_addr_11 <= _GEN_622;
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_2) begin // @[Conditional.scala 39:67]
        L1_wrEna_0 <= _GEN_56;
      end else if (_T_13) begin // @[Conditional.scala 39:67]
        if (count == 10'h34) begin // @[FSM.scala 276:27]
          L1_wrEna_0 <= 1'h0; // @[FSM.scala 278:23]
        end else begin
          L1_wrEna_0 <= _GEN_206;
        end
      end else if (_T_32) begin // @[Conditional.scala 39:67]
        L1_wrEna_0 <= _GEN_623;
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_2) begin // @[Conditional.scala 39:67]
        L1_wrEna_1 <= _GEN_58;
      end else if (_T_13) begin // @[Conditional.scala 39:67]
        if (count == 10'h34) begin // @[FSM.scala 276:27]
          L1_wrEna_1 <= 1'h0; // @[FSM.scala 278:23]
        end else begin
          L1_wrEna_1 <= _GEN_208;
        end
      end else if (_T_32) begin // @[Conditional.scala 39:67]
        L1_wrEna_1 <= _GEN_624;
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_2) begin // @[Conditional.scala 39:67]
        L1_wrEna_2 <= _GEN_60;
      end else if (_T_13) begin // @[Conditional.scala 39:67]
        if (count == 10'h34) begin // @[FSM.scala 276:27]
          L1_wrEna_2 <= 1'h0; // @[FSM.scala 278:23]
        end else begin
          L1_wrEna_2 <= _GEN_209;
        end
      end else if (_T_32) begin // @[Conditional.scala 39:67]
        L1_wrEna_2 <= _GEN_625;
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_2) begin // @[Conditional.scala 39:67]
        L1_wrEna_3 <= _GEN_62;
      end else if (_T_13) begin // @[Conditional.scala 39:67]
        if (count == 10'h34) begin // @[FSM.scala 276:27]
          L1_wrEna_3 <= 1'h0; // @[FSM.scala 278:23]
        end else begin
          L1_wrEna_3 <= _GEN_210;
        end
      end else if (_T_32) begin // @[Conditional.scala 39:67]
        L1_wrEna_3 <= _GEN_626;
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_2) begin // @[Conditional.scala 39:67]
        L1_wrEna_4 <= _GEN_64;
      end else if (_T_13) begin // @[Conditional.scala 39:67]
        if (count == 10'h34) begin // @[FSM.scala 276:27]
          L1_wrEna_4 <= 1'h0; // @[FSM.scala 278:23]
        end else begin
          L1_wrEna_4 <= _GEN_211;
        end
      end else if (_T_32) begin // @[Conditional.scala 39:67]
        L1_wrEna_4 <= _GEN_627;
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_2) begin // @[Conditional.scala 39:67]
        L1_wrEna_5 <= _GEN_66;
      end else if (_T_13) begin // @[Conditional.scala 39:67]
        if (count == 10'h34) begin // @[FSM.scala 276:27]
          L1_wrEna_5 <= 1'h0; // @[FSM.scala 278:23]
        end else begin
          L1_wrEna_5 <= _GEN_212;
        end
      end else if (_T_32) begin // @[Conditional.scala 39:67]
        L1_wrEna_5 <= _GEN_628;
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_2) begin // @[Conditional.scala 39:67]
        L1_wrEna_6 <= _GEN_68;
      end else if (_T_13) begin // @[Conditional.scala 39:67]
        if (count == 10'h34) begin // @[FSM.scala 276:27]
          L1_wrEna_6 <= 1'h0; // @[FSM.scala 278:23]
        end else begin
          L1_wrEna_6 <= _GEN_213;
        end
      end else if (_T_32) begin // @[Conditional.scala 39:67]
        L1_wrEna_6 <= _GEN_629;
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_2) begin // @[Conditional.scala 39:67]
        L1_wrEna_7 <= _GEN_70;
      end else if (_T_13) begin // @[Conditional.scala 39:67]
        if (count == 10'h34) begin // @[FSM.scala 276:27]
          L1_wrEna_7 <= 1'h0; // @[FSM.scala 278:23]
        end else begin
          L1_wrEna_7 <= _GEN_214;
        end
      end else if (_T_32) begin // @[Conditional.scala 39:67]
        L1_wrEna_7 <= _GEN_630;
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_2) begin // @[Conditional.scala 39:67]
        L1_wrEna_8 <= _GEN_72;
      end else if (_T_13) begin // @[Conditional.scala 39:67]
        if (count == 10'h34) begin // @[FSM.scala 276:27]
          L1_wrEna_8 <= 1'h0; // @[FSM.scala 278:23]
        end else begin
          L1_wrEna_8 <= _GEN_215;
        end
      end else if (_T_32) begin // @[Conditional.scala 39:67]
        L1_wrEna_8 <= _GEN_631;
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_2) begin // @[Conditional.scala 39:67]
        L1_wrEna_9 <= _GEN_74;
      end else if (_T_13) begin // @[Conditional.scala 39:67]
        if (count == 10'h34) begin // @[FSM.scala 276:27]
          L1_wrEna_9 <= 1'h0; // @[FSM.scala 278:23]
        end else begin
          L1_wrEna_9 <= _GEN_216;
        end
      end else if (_T_32) begin // @[Conditional.scala 39:67]
        L1_wrEna_9 <= _GEN_632;
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_2) begin // @[Conditional.scala 39:67]
        L1_wrEna_10 <= _GEN_76;
      end else if (_T_13) begin // @[Conditional.scala 39:67]
        if (count == 10'h34) begin // @[FSM.scala 276:27]
          L1_wrEna_10 <= 1'h0; // @[FSM.scala 278:23]
        end else begin
          L1_wrEna_10 <= _GEN_217;
        end
      end else if (_T_32) begin // @[Conditional.scala 39:67]
        L1_wrEna_10 <= _GEN_633;
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_2) begin // @[Conditional.scala 39:67]
        L1_wrEna_11 <= _GEN_78;
      end else if (_T_13) begin // @[Conditional.scala 39:67]
        if (count == 10'h34) begin // @[FSM.scala 276:27]
          L1_wrEna_11 <= 1'h0; // @[FSM.scala 278:23]
        end else begin
          L1_wrEna_11 <= _GEN_218;
        end
      end else if (_T_32) begin // @[Conditional.scala 39:67]
        L1_wrEna_11 <= _GEN_634;
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          if (_T_5) begin // @[FSM.scala 235:26]
            PEArray_ctrl_0_mask <= 12'h0; // @[FSM.scala 237:32]
          end else begin
            PEArray_ctrl_0_mask <= _GEN_87;
          end
        end else if (_T_32) begin // @[Conditional.scala 39:67]
          PEArray_ctrl_0_mask <= _GEN_291;
        end else begin
          PEArray_ctrl_0_mask <= _GEN_2035;
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          if (_T_5) begin // @[FSM.scala 235:26]
            PEArray_ctrl_1_mask <= 12'h0; // @[FSM.scala 237:32]
          end else begin
            PEArray_ctrl_1_mask <= _GEN_89;
          end
        end else if (_T_32) begin // @[Conditional.scala 39:67]
          PEArray_ctrl_1_mask <= _GEN_292;
        end else begin
          PEArray_ctrl_1_mask <= _GEN_2036;
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          if (_T_3) begin // @[FSM.scala 223:26]
            PEArray_ctrl_2_control <= 3'h1; // @[FSM.scala 225:35]
          end
        end else if (_T_32) begin // @[Conditional.scala 39:67]
          PEArray_ctrl_2_control <= _GEN_289;
        end else begin
          PEArray_ctrl_2_control <= _GEN_2029;
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_13)) begin // @[Conditional.scala 39:67]
          if (!(_T_32)) begin // @[Conditional.scala 39:67]
            PEArray_ctrl_2_count <= _GEN_2031;
          end
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_13)) begin // @[Conditional.scala 39:67]
          if (!(_T_32)) begin // @[Conditional.scala 39:67]
            PEArray_ctrl_2_L0index <= _GEN_2032;
          end
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          if (_T_5) begin // @[FSM.scala 235:26]
            PEArray_ctrl_2_mask <= 12'h0; // @[FSM.scala 237:32]
          end else begin
            PEArray_ctrl_2_mask <= _GEN_91;
          end
        end else if (_T_32) begin // @[Conditional.scala 39:67]
          PEArray_ctrl_2_mask <= _GEN_293;
        end else begin
          PEArray_ctrl_2_mask <= _GEN_2030;
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_13)) begin // @[Conditional.scala 39:67]
          if (!(_T_32)) begin // @[Conditional.scala 39:67]
            PEArray_ctrl_2_gru_out_width <= _GEN_2052;
          end
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          if (count == 10'h4) begin // @[FSM.scala 247:26]
            BNArray_ctrl_0 <= 2'h0; // @[FSM.scala 251:27]
          end
        end else if (_T_32) begin // @[Conditional.scala 39:67]
          BNArray_ctrl_0 <= _GEN_254;
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          if (count == 10'h4) begin // @[FSM.scala 247:26]
            BNArray_ctrl_1 <= 2'h0; // @[FSM.scala 251:27]
          end
        end else if (_T_32) begin // @[Conditional.scala 39:67]
          BNArray_ctrl_1 <= _GEN_257;
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          if (count == 10'h4) begin // @[FSM.scala 247:26]
            BNArray_ctrl_2 <= 2'h0; // @[FSM.scala 251:27]
          end
        end else if (_T_32) begin // @[Conditional.scala 39:67]
          BNArray_ctrl_2 <= _GEN_260;
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          if (count == 10'h4) begin // @[FSM.scala 247:26]
            BNArray_ctrl_3 <= 2'h0; // @[FSM.scala 251:27]
          end
        end else if (_T_32) begin // @[Conditional.scala 39:67]
          BNArray_ctrl_3 <= _GEN_263;
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          if (count == 10'h4) begin // @[FSM.scala 247:26]
            BNArray_ctrl_4 <= 2'h0; // @[FSM.scala 251:27]
          end
        end else if (_T_32) begin // @[Conditional.scala 39:67]
          BNArray_ctrl_4 <= _GEN_266;
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          if (count == 10'h4) begin // @[FSM.scala 247:26]
            BNArray_ctrl_5 <= 2'h0; // @[FSM.scala 251:27]
          end
        end else if (_T_32) begin // @[Conditional.scala 39:67]
          BNArray_ctrl_5 <= _GEN_269;
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          if (count == 10'h4) begin // @[FSM.scala 247:26]
            BNArray_ctrl_6 <= 2'h0; // @[FSM.scala 251:27]
          end
        end else if (_T_32) begin // @[Conditional.scala 39:67]
          BNArray_ctrl_6 <= _GEN_272;
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          if (count == 10'h4) begin // @[FSM.scala 247:26]
            BNArray_ctrl_7 <= 2'h0; // @[FSM.scala 251:27]
          end
        end else if (_T_32) begin // @[Conditional.scala 39:67]
          BNArray_ctrl_7 <= _GEN_275;
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          if (count == 10'h4) begin // @[FSM.scala 247:26]
            BNArray_ctrl_8 <= 2'h0; // @[FSM.scala 251:27]
          end
        end else if (_T_32) begin // @[Conditional.scala 39:67]
          BNArray_ctrl_8 <= _GEN_278;
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          if (count == 10'h4) begin // @[FSM.scala 247:26]
            BNArray_ctrl_9 <= 2'h0; // @[FSM.scala 251:27]
          end
        end else if (_T_32) begin // @[Conditional.scala 39:67]
          BNArray_ctrl_9 <= _GEN_281;
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          if (count == 10'h4) begin // @[FSM.scala 247:26]
            BNArray_ctrl_10 <= 2'h0; // @[FSM.scala 251:27]
          end
        end else if (_T_32) begin // @[Conditional.scala 39:67]
          BNArray_ctrl_10 <= _GEN_284;
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          if (count == 10'h4) begin // @[FSM.scala 247:26]
            BNArray_ctrl_11 <= 2'h0; // @[FSM.scala 251:27]
          end
        end else if (_T_32) begin // @[Conditional.scala 39:67]
          BNArray_ctrl_11 <= _GEN_287;
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_13)) begin // @[Conditional.scala 39:67]
          if (!(_T_32)) begin // @[Conditional.scala 39:67]
            BN_Unit_ctrl <= _GEN_2054;
          end
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          if (count == 10'h4) begin // @[FSM.scala 247:26]
            Relu6Array_ctrl_0 <= 1'h0; // @[FSM.scala 252:30]
          end
        end else if (_T_32) begin // @[Conditional.scala 39:67]
          Relu6Array_ctrl_0 <= _GEN_255;
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          if (count == 10'h4) begin // @[FSM.scala 247:26]
            Relu6Array_ctrl_1 <= 1'h0; // @[FSM.scala 252:30]
          end
        end else if (_T_32) begin // @[Conditional.scala 39:67]
          Relu6Array_ctrl_1 <= _GEN_258;
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          if (count == 10'h4) begin // @[FSM.scala 247:26]
            Relu6Array_ctrl_2 <= 1'h0; // @[FSM.scala 252:30]
          end
        end else if (_T_32) begin // @[Conditional.scala 39:67]
          Relu6Array_ctrl_2 <= _GEN_261;
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          if (count == 10'h4) begin // @[FSM.scala 247:26]
            Relu6Array_ctrl_3 <= 1'h0; // @[FSM.scala 252:30]
          end
        end else if (_T_32) begin // @[Conditional.scala 39:67]
          Relu6Array_ctrl_3 <= _GEN_264;
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          if (count == 10'h4) begin // @[FSM.scala 247:26]
            Relu6Array_ctrl_4 <= 1'h0; // @[FSM.scala 252:30]
          end
        end else if (_T_32) begin // @[Conditional.scala 39:67]
          Relu6Array_ctrl_4 <= _GEN_267;
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          if (count == 10'h4) begin // @[FSM.scala 247:26]
            Relu6Array_ctrl_5 <= 1'h0; // @[FSM.scala 252:30]
          end
        end else if (_T_32) begin // @[Conditional.scala 39:67]
          Relu6Array_ctrl_5 <= _GEN_270;
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          if (count == 10'h4) begin // @[FSM.scala 247:26]
            Relu6Array_ctrl_6 <= 1'h0; // @[FSM.scala 252:30]
          end
        end else if (_T_32) begin // @[Conditional.scala 39:67]
          Relu6Array_ctrl_6 <= _GEN_273;
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          if (count == 10'h4) begin // @[FSM.scala 247:26]
            Relu6Array_ctrl_7 <= 1'h0; // @[FSM.scala 252:30]
          end
        end else if (_T_32) begin // @[Conditional.scala 39:67]
          Relu6Array_ctrl_7 <= _GEN_276;
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          if (count == 10'h4) begin // @[FSM.scala 247:26]
            Relu6Array_ctrl_8 <= 1'h0; // @[FSM.scala 252:30]
          end
        end else if (_T_32) begin // @[Conditional.scala 39:67]
          Relu6Array_ctrl_8 <= _GEN_279;
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          if (count == 10'h4) begin // @[FSM.scala 247:26]
            Relu6Array_ctrl_9 <= 1'h0; // @[FSM.scala 252:30]
          end
        end else if (_T_32) begin // @[Conditional.scala 39:67]
          Relu6Array_ctrl_9 <= _GEN_282;
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          if (count == 10'h4) begin // @[FSM.scala 247:26]
            Relu6Array_ctrl_10 <= 1'h0; // @[FSM.scala 252:30]
          end
        end else if (_T_32) begin // @[Conditional.scala 39:67]
          Relu6Array_ctrl_10 <= _GEN_285;
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          if (count == 10'h4) begin // @[FSM.scala 247:26]
            Relu6Array_ctrl_11 <= 1'h0; // @[FSM.scala 252:30]
          end
        end else if (_T_32) begin // @[Conditional.scala 39:67]
          Relu6Array_ctrl_11 <= _GEN_288;
        end
      end
    end
    if (reset) begin // @[FSM.scala 74:35]
      PE_above_data_ctrl <= 2'h0; // @[FSM.scala 74:35]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          PE_above_data_ctrl <= _GEN_104;
        end else begin
          PE_above_data_ctrl <= _GEN_2093;
        end
      end
    end
    if (reset) begin // @[FSM.scala 75:32]
      Activation_ctrl <= 2'h0; // @[FSM.scala 75:32]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_13)) begin // @[Conditional.scala 39:67]
          Activation_ctrl <= _GEN_2155;
        end
      end
    end
    if (reset) begin // @[FSM.scala 77:36]
      Ht_to_PE_control <= 3'h0; // @[FSM.scala 77:36]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_13)) begin // @[Conditional.scala 39:67]
          Ht_to_PE_control <= _GEN_2150;
        end
      end
    end
    if (reset) begin // @[FSM.scala 79:36]
      Ht_wrEna <= 1'h0; // @[FSM.scala 79:36]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_13)) begin // @[Conditional.scala 39:67]
          Ht_wrEna <= _GEN_2168;
        end
      end
    end
    if (reset) begin // @[FSM.scala 80:36]
      Ht_wrAddr <= 6'h0; // @[FSM.scala 80:36]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_13)) begin // @[Conditional.scala 39:67]
          Ht_wrAddr <= _GEN_2167;
        end
      end
    end
    if (reset) begin // @[FSM.scala 81:36]
      Zt_rdAddr <= 6'h0; // @[FSM.scala 81:36]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_13)) begin // @[Conditional.scala 39:67]
          Zt_rdAddr <= _GEN_2163;
        end
      end
    end
    if (reset) begin // @[FSM.scala 82:36]
      Zt_wrEna <= 1'h0; // @[FSM.scala 82:36]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_13)) begin // @[Conditional.scala 39:67]
          Zt_wrEna <= _GEN_2156;
        end
      end
    end
    if (reset) begin // @[FSM.scala 83:36]
      Zt_wrAddr <= 6'h0; // @[FSM.scala 83:36]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_13)) begin // @[Conditional.scala 39:67]
          Zt_wrAddr <= _GEN_2153;
        end
      end
    end
    if (reset) begin // @[FSM.scala 84:36]
      Rt_rdAddr <= 6'h0; // @[FSM.scala 84:36]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_13)) begin // @[Conditional.scala 39:67]
          Rt_rdAddr <= _GEN_2164;
        end
      end
    end
    if (reset) begin // @[FSM.scala 85:36]
      Rt_wrEna <= 1'h0; // @[FSM.scala 85:36]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_13)) begin // @[Conditional.scala 39:67]
          Rt_wrEna <= _GEN_2158;
        end
      end
    end
    if (reset) begin // @[FSM.scala 86:36]
      Rt_wrAddr <= 6'h0; // @[FSM.scala 86:36]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_13)) begin // @[Conditional.scala 39:67]
          Rt_wrAddr <= _GEN_2157;
        end
      end
    end
    if (reset) begin // @[FSM.scala 87:36]
      WhXt_rdAddr <= 6'h0; // @[FSM.scala 87:36]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_13)) begin // @[Conditional.scala 39:67]
          WhXt_rdAddr <= _GEN_2165;
        end
      end
    end
    if (reset) begin // @[FSM.scala 88:36]
      WhXt_wrEna <= 1'h0; // @[FSM.scala 88:36]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_13)) begin // @[Conditional.scala 39:67]
          WhXt_wrEna <= _GEN_2160;
        end
      end
    end
    if (reset) begin // @[FSM.scala 89:36]
      WhXt_wrAddr <= 6'h0; // @[FSM.scala 89:36]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_13)) begin // @[Conditional.scala 39:67]
          WhXt_wrAddr <= _GEN_2159;
        end
      end
    end
    if (reset) begin // @[FSM.scala 90:36]
      Uhht_1_rdAddr <= 6'h0; // @[FSM.scala 90:36]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_13)) begin // @[Conditional.scala 39:67]
          Uhht_1_rdAddr <= _GEN_2166;
        end
      end
    end
    if (reset) begin // @[FSM.scala 91:36]
      Uhht_1_wrEna <= 1'h0; // @[FSM.scala 91:36]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_13)) begin // @[Conditional.scala 39:67]
          Uhht_1_wrEna <= _GEN_2162;
        end
      end
    end
    if (reset) begin // @[FSM.scala 92:36]
      Uhht_1_wrAddr <= 6'h0; // @[FSM.scala 92:36]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_13)) begin // @[Conditional.scala 39:67]
          Uhht_1_wrAddr <= _GEN_2161;
        end
      end
    end
    if (reset) begin // @[FSM.scala 94:38]
      FC_temp_to_PE_control <= 3'h0; // @[FSM.scala 94:38]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_13)) begin // @[Conditional.scala 39:67]
          FC_temp_to_PE_control <= _GEN_2173;
        end
      end
    end
    if (reset) begin // @[FSM.scala 96:38]
      FC_temp_wrEna <= 1'h0; // @[FSM.scala 96:38]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_13)) begin // @[Conditional.scala 39:67]
          FC_temp_wrEna <= _GEN_2172;
        end
      end
    end
    if (reset) begin // @[FSM.scala 97:38]
      FC_temp_wrAddr <= 6'h0; // @[FSM.scala 97:38]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_13)) begin // @[Conditional.scala 39:67]
          FC_temp_wrAddr <= _GEN_2171;
        end
      end
    end
    if (reset) begin // @[FSM.scala 99:38]
      Result_wrEna <= 1'h0; // @[FSM.scala 99:38]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_13)) begin // @[Conditional.scala 39:67]
          Result_wrEna <= _GEN_2175;
        end
      end
    end
    if (reset) begin // @[FSM.scala 100:38]
      Result_wrAddr <= 4'h0; // @[FSM.scala 100:38]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_13)) begin // @[Conditional.scala 39:67]
          Result_wrAddr <= _GEN_2174;
        end
      end
    end
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_2) begin // @[Conditional.scala 39:67]
        if (io_Input_Valid & io_Input_Ready) begin // @[FSM.scala 202:67]
          Data_temp <= io_Input_Data; // @[FSM.scala 203:19]
        end
      end
    end
    Data_temp_used <= reset | _GEN_2386; // @[FSM.scala 105:31 FSM.scala 105:31]
    if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_2) begin // @[Conditional.scala 39:67]
        if (~Data_temp_used) begin // @[FSM.scala 179:39]
          if (count >= 10'h2 & count <= 10'hf) begin // @[FSM.scala 189:44]
            L1_wr_data <= Data_temp; // @[FSM.scala 190:22]
          end else begin
            L1_wr_data <= _GEN_3;
          end
        end
      end
    end
    if (reset) begin // @[FSM.scala 159:22]
      state <= 3'h0; // @[FSM.scala 159:22]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_Start) begin // @[FSM.scala 170:32]
        state <= 3'h1; // @[FSM.scala 171:15]
      end
    end else if (_T_2) begin // @[Conditional.scala 39:67]
      if (count == 10'h10) begin // @[FSM.scala 207:27]
        state <= 3'h2; // @[FSM.scala 208:15]
      end
    end else if (_T_13) begin // @[Conditional.scala 39:67]
      state <= _GEN_233;
    end else begin
      state <= _GEN_2147;
    end
    if (reset) begin // @[FSM.scala 160:26]
      gru_state <= 4'h0; // @[FSM.scala 160:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_13)) begin // @[Conditional.scala 39:67]
          gru_state <= _GEN_2151;
        end
      end
    end
    if (reset) begin // @[FSM.scala 161:22]
      count <= 10'h0; // @[FSM.scala 161:22]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_2) begin // @[Conditional.scala 39:67]
        if (io_Input_Valid & io_Input_Ready) begin // @[FSM.scala 202:67]
          count <= _count_T_1; // @[FSM.scala 205:15]
        end
      end else if (_T_13) begin // @[Conditional.scala 39:67]
        count <= _GEN_231;
      end else begin
        count <= _GEN_2077;
      end
    end
    if (reset) begin // @[FSM.scala 162:23]
      count1 <= 7'h0; // @[FSM.scala 162:23]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[Conditional.scala 39:67]
          count1 <= _GEN_232;
        end else begin
          count1 <= _GEN_2078;
        end
      end
    end
    if (reset) begin // @[FSM.scala 164:26]
      gru_count <= 6'h0; // @[FSM.scala 164:26]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_13)) begin // @[Conditional.scala 39:67]
          gru_count <= _GEN_2169;
        end
      end
    end
    if (reset) begin // @[FSM.scala 165:27]
      read_index <= 4'h0; // @[FSM.scala 165:27]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_13)) begin // @[Conditional.scala 39:67]
          read_index <= _GEN_2133;
        end
      end
    end
    if (reset) begin // @[FSM.scala 166:25]
      fc_state <= 2'h0; // @[FSM.scala 166:25]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (!(_T_2)) begin // @[Conditional.scala 39:67]
        if (!(_T_13)) begin // @[Conditional.scala 39:67]
          fc_state <= _GEN_2170;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  L1_rd_addr_0 = _RAND_0[11:0];
  _RAND_1 = {1{`RANDOM}};
  L1_rd_addr_1 = _RAND_1[11:0];
  _RAND_2 = {1{`RANDOM}};
  L1_rd_addr_2 = _RAND_2[11:0];
  _RAND_3 = {1{`RANDOM}};
  L1_rd_addr_3 = _RAND_3[11:0];
  _RAND_4 = {1{`RANDOM}};
  L1_rd_addr_4 = _RAND_4[11:0];
  _RAND_5 = {1{`RANDOM}};
  L1_rd_addr_5 = _RAND_5[11:0];
  _RAND_6 = {1{`RANDOM}};
  L1_rd_addr_6 = _RAND_6[11:0];
  _RAND_7 = {1{`RANDOM}};
  L1_rd_addr_7 = _RAND_7[11:0];
  _RAND_8 = {1{`RANDOM}};
  L1_rd_addr_8 = _RAND_8[11:0];
  _RAND_9 = {1{`RANDOM}};
  L1_rd_addr_9 = _RAND_9[11:0];
  _RAND_10 = {1{`RANDOM}};
  L1_rd_addr_10 = _RAND_10[11:0];
  _RAND_11 = {1{`RANDOM}};
  L1_rd_addr_11 = _RAND_11[11:0];
  _RAND_12 = {1{`RANDOM}};
  PE_rd_data_mux = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  L1_wr_addr_0 = _RAND_13[11:0];
  _RAND_14 = {1{`RANDOM}};
  L1_wr_addr_1 = _RAND_14[11:0];
  _RAND_15 = {1{`RANDOM}};
  L1_wr_addr_2 = _RAND_15[11:0];
  _RAND_16 = {1{`RANDOM}};
  L1_wr_addr_3 = _RAND_16[11:0];
  _RAND_17 = {1{`RANDOM}};
  L1_wr_addr_4 = _RAND_17[11:0];
  _RAND_18 = {1{`RANDOM}};
  L1_wr_addr_5 = _RAND_18[11:0];
  _RAND_19 = {1{`RANDOM}};
  L1_wr_addr_6 = _RAND_19[11:0];
  _RAND_20 = {1{`RANDOM}};
  L1_wr_addr_7 = _RAND_20[11:0];
  _RAND_21 = {1{`RANDOM}};
  L1_wr_addr_8 = _RAND_21[11:0];
  _RAND_22 = {1{`RANDOM}};
  L1_wr_addr_9 = _RAND_22[11:0];
  _RAND_23 = {1{`RANDOM}};
  L1_wr_addr_10 = _RAND_23[11:0];
  _RAND_24 = {1{`RANDOM}};
  L1_wr_addr_11 = _RAND_24[11:0];
  _RAND_25 = {1{`RANDOM}};
  L1_wrEna_0 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  L1_wrEna_1 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  L1_wrEna_2 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  L1_wrEna_3 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  L1_wrEna_4 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  L1_wrEna_5 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  L1_wrEna_6 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  L1_wrEna_7 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  L1_wrEna_8 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  L1_wrEna_9 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  L1_wrEna_10 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  L1_wrEna_11 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  PEArray_ctrl_0_mask = _RAND_37[11:0];
  _RAND_38 = {1{`RANDOM}};
  PEArray_ctrl_1_mask = _RAND_38[11:0];
  _RAND_39 = {1{`RANDOM}};
  PEArray_ctrl_2_control = _RAND_39[2:0];
  _RAND_40 = {1{`RANDOM}};
  PEArray_ctrl_2_count = _RAND_40[9:0];
  _RAND_41 = {1{`RANDOM}};
  PEArray_ctrl_2_L0index = _RAND_41[5:0];
  _RAND_42 = {1{`RANDOM}};
  PEArray_ctrl_2_mask = _RAND_42[11:0];
  _RAND_43 = {1{`RANDOM}};
  PEArray_ctrl_2_gru_out_width = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  BNArray_ctrl_0 = _RAND_44[1:0];
  _RAND_45 = {1{`RANDOM}};
  BNArray_ctrl_1 = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  BNArray_ctrl_2 = _RAND_46[1:0];
  _RAND_47 = {1{`RANDOM}};
  BNArray_ctrl_3 = _RAND_47[1:0];
  _RAND_48 = {1{`RANDOM}};
  BNArray_ctrl_4 = _RAND_48[1:0];
  _RAND_49 = {1{`RANDOM}};
  BNArray_ctrl_5 = _RAND_49[1:0];
  _RAND_50 = {1{`RANDOM}};
  BNArray_ctrl_6 = _RAND_50[1:0];
  _RAND_51 = {1{`RANDOM}};
  BNArray_ctrl_7 = _RAND_51[1:0];
  _RAND_52 = {1{`RANDOM}};
  BNArray_ctrl_8 = _RAND_52[1:0];
  _RAND_53 = {1{`RANDOM}};
  BNArray_ctrl_9 = _RAND_53[1:0];
  _RAND_54 = {1{`RANDOM}};
  BNArray_ctrl_10 = _RAND_54[1:0];
  _RAND_55 = {1{`RANDOM}};
  BNArray_ctrl_11 = _RAND_55[1:0];
  _RAND_56 = {1{`RANDOM}};
  BN_Unit_ctrl = _RAND_56[1:0];
  _RAND_57 = {1{`RANDOM}};
  Relu6Array_ctrl_0 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  Relu6Array_ctrl_1 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  Relu6Array_ctrl_2 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  Relu6Array_ctrl_3 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  Relu6Array_ctrl_4 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  Relu6Array_ctrl_5 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  Relu6Array_ctrl_6 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  Relu6Array_ctrl_7 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  Relu6Array_ctrl_8 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  Relu6Array_ctrl_9 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  Relu6Array_ctrl_10 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  Relu6Array_ctrl_11 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  PE_above_data_ctrl = _RAND_69[1:0];
  _RAND_70 = {1{`RANDOM}};
  Activation_ctrl = _RAND_70[1:0];
  _RAND_71 = {1{`RANDOM}};
  Ht_to_PE_control = _RAND_71[2:0];
  _RAND_72 = {1{`RANDOM}};
  Ht_wrEna = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  Ht_wrAddr = _RAND_73[5:0];
  _RAND_74 = {1{`RANDOM}};
  Zt_rdAddr = _RAND_74[5:0];
  _RAND_75 = {1{`RANDOM}};
  Zt_wrEna = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  Zt_wrAddr = _RAND_76[5:0];
  _RAND_77 = {1{`RANDOM}};
  Rt_rdAddr = _RAND_77[5:0];
  _RAND_78 = {1{`RANDOM}};
  Rt_wrEna = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  Rt_wrAddr = _RAND_79[5:0];
  _RAND_80 = {1{`RANDOM}};
  WhXt_rdAddr = _RAND_80[5:0];
  _RAND_81 = {1{`RANDOM}};
  WhXt_wrEna = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  WhXt_wrAddr = _RAND_82[5:0];
  _RAND_83 = {1{`RANDOM}};
  Uhht_1_rdAddr = _RAND_83[5:0];
  _RAND_84 = {1{`RANDOM}};
  Uhht_1_wrEna = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  Uhht_1_wrAddr = _RAND_85[5:0];
  _RAND_86 = {1{`RANDOM}};
  FC_temp_to_PE_control = _RAND_86[2:0];
  _RAND_87 = {1{`RANDOM}};
  FC_temp_wrEna = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  FC_temp_wrAddr = _RAND_88[5:0];
  _RAND_89 = {1{`RANDOM}};
  Result_wrEna = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  Result_wrAddr = _RAND_90[3:0];
  _RAND_91 = {1{`RANDOM}};
  Data_temp = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  Data_temp_used = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  L1_wr_data = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  state = _RAND_94[2:0];
  _RAND_95 = {1{`RANDOM}};
  gru_state = _RAND_95[3:0];
  _RAND_96 = {1{`RANDOM}};
  count = _RAND_96[9:0];
  _RAND_97 = {1{`RANDOM}};
  count1 = _RAND_97[6:0];
  _RAND_98 = {1{`RANDOM}};
  gru_count = _RAND_98[5:0];
  _RAND_99 = {1{`RANDOM}};
  read_index = _RAND_99[3:0];
  _RAND_100 = {1{`RANDOM}};
  fc_state = _RAND_100[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BN_Unit(
  input         clock,
  input         reset,
  input  [15:0] io_input,
  input  [1:0]  io_control,
  output [15:0] io_output
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] FP16MAC_io_a; // @[Unit.scala 21:23]
  wire [15:0] FP16MAC_io_b; // @[Unit.scala 21:23]
  wire [15:0] FP16MAC_io_c; // @[Unit.scala 21:23]
  wire [15:0] FP16MAC_io_out; // @[Unit.scala 21:23]
  reg [15:0] output_reg; // @[Unit.scala 17:27]
  wire [15:0] _GEN_9 = FP16MAC_io_out; // @[Unit.scala 43:32 Unit.scala 47:16 Unit.scala 53:16]
  wire [13:0] _GEN_15 = io_control == 2'h0 ? 14'h0 : 14'h3c00; // @[Unit.scala 31:27 Unit.scala 33:18]
  FP16MulAdder FP16MAC ( // @[Unit.scala 21:23]
    .io_a(FP16MAC_io_a),
    .io_b(FP16MAC_io_b),
    .io_c(FP16MAC_io_c),
    .io_out(FP16MAC_io_out)
  );
  assign io_output = output_reg; // @[Unit.scala 18:13]
  assign FP16MAC_io_a = io_control == 2'h0 ? 16'h0 : io_input; // @[Unit.scala 31:27 Unit.scala 32:18]
  assign FP16MAC_io_b = {{2'd0}, _GEN_15}; // @[Unit.scala 31:27 Unit.scala 33:18]
  assign FP16MAC_io_c = 16'h0; // @[Unit.scala 31:27 Unit.scala 34:18]
  always @(posedge clock) begin
    if (reset) begin // @[Unit.scala 17:27]
      output_reg <= 16'h0; // @[Unit.scala 17:27]
    end else if (io_control == 2'h0) begin // @[Unit.scala 31:27]
      output_reg <= io_input; // @[Unit.scala 35:16]
    end else if (io_control == 2'h1) begin // @[Unit.scala 37:32]
      output_reg <= FP16MAC_io_out; // @[Unit.scala 41:16]
    end else begin
      output_reg <= _GEN_9;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  output_reg = _RAND_0[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BN_Unit_Array(
  input         clock,
  input         reset,
  input  [15:0] io_from_PE_0,
  input  [15:0] io_from_PE_1,
  input  [15:0] io_from_PE_2,
  input  [15:0] io_from_PE_3,
  input  [15:0] io_from_PE_4,
  input  [15:0] io_from_PE_5,
  input  [15:0] io_from_PE_6,
  input  [15:0] io_from_PE_7,
  input  [15:0] io_from_PE_8,
  input  [15:0] io_from_PE_9,
  input  [15:0] io_from_PE_10,
  input  [15:0] io_from_PE_11,
  input  [1:0]  io_control_0,
  input  [1:0]  io_control_1,
  input  [1:0]  io_control_2,
  input  [1:0]  io_control_3,
  input  [1:0]  io_control_4,
  input  [1:0]  io_control_5,
  input  [1:0]  io_control_6,
  input  [1:0]  io_control_7,
  input  [1:0]  io_control_8,
  input  [1:0]  io_control_9,
  input  [1:0]  io_control_10,
  input  [1:0]  io_control_11,
  output [15:0] io_to_Relu6_0,
  output [15:0] io_to_Relu6_1,
  output [15:0] io_to_Relu6_2,
  output [15:0] io_to_Relu6_3,
  output [15:0] io_to_Relu6_4,
  output [15:0] io_to_Relu6_5,
  output [15:0] io_to_Relu6_6,
  output [15:0] io_to_Relu6_7,
  output [15:0] io_to_Relu6_8,
  output [15:0] io_to_Relu6_9,
  output [15:0] io_to_Relu6_10,
  output [15:0] io_to_Relu6_11
);
  wire  BN_Array_0_clock; // @[Unit.scala 68:37]
  wire  BN_Array_0_reset; // @[Unit.scala 68:37]
  wire [15:0] BN_Array_0_io_input; // @[Unit.scala 68:37]
  wire [1:0] BN_Array_0_io_control; // @[Unit.scala 68:37]
  wire [15:0] BN_Array_0_io_output; // @[Unit.scala 68:37]
  wire  BN_Array_1_clock; // @[Unit.scala 68:37]
  wire  BN_Array_1_reset; // @[Unit.scala 68:37]
  wire [15:0] BN_Array_1_io_input; // @[Unit.scala 68:37]
  wire [1:0] BN_Array_1_io_control; // @[Unit.scala 68:37]
  wire [15:0] BN_Array_1_io_output; // @[Unit.scala 68:37]
  wire  BN_Array_2_clock; // @[Unit.scala 68:37]
  wire  BN_Array_2_reset; // @[Unit.scala 68:37]
  wire [15:0] BN_Array_2_io_input; // @[Unit.scala 68:37]
  wire [1:0] BN_Array_2_io_control; // @[Unit.scala 68:37]
  wire [15:0] BN_Array_2_io_output; // @[Unit.scala 68:37]
  wire  BN_Array_3_clock; // @[Unit.scala 68:37]
  wire  BN_Array_3_reset; // @[Unit.scala 68:37]
  wire [15:0] BN_Array_3_io_input; // @[Unit.scala 68:37]
  wire [1:0] BN_Array_3_io_control; // @[Unit.scala 68:37]
  wire [15:0] BN_Array_3_io_output; // @[Unit.scala 68:37]
  wire  BN_Array_4_clock; // @[Unit.scala 68:37]
  wire  BN_Array_4_reset; // @[Unit.scala 68:37]
  wire [15:0] BN_Array_4_io_input; // @[Unit.scala 68:37]
  wire [1:0] BN_Array_4_io_control; // @[Unit.scala 68:37]
  wire [15:0] BN_Array_4_io_output; // @[Unit.scala 68:37]
  wire  BN_Array_5_clock; // @[Unit.scala 68:37]
  wire  BN_Array_5_reset; // @[Unit.scala 68:37]
  wire [15:0] BN_Array_5_io_input; // @[Unit.scala 68:37]
  wire [1:0] BN_Array_5_io_control; // @[Unit.scala 68:37]
  wire [15:0] BN_Array_5_io_output; // @[Unit.scala 68:37]
  wire  BN_Array_6_clock; // @[Unit.scala 68:37]
  wire  BN_Array_6_reset; // @[Unit.scala 68:37]
  wire [15:0] BN_Array_6_io_input; // @[Unit.scala 68:37]
  wire [1:0] BN_Array_6_io_control; // @[Unit.scala 68:37]
  wire [15:0] BN_Array_6_io_output; // @[Unit.scala 68:37]
  wire  BN_Array_7_clock; // @[Unit.scala 68:37]
  wire  BN_Array_7_reset; // @[Unit.scala 68:37]
  wire [15:0] BN_Array_7_io_input; // @[Unit.scala 68:37]
  wire [1:0] BN_Array_7_io_control; // @[Unit.scala 68:37]
  wire [15:0] BN_Array_7_io_output; // @[Unit.scala 68:37]
  wire  BN_Array_8_clock; // @[Unit.scala 68:37]
  wire  BN_Array_8_reset; // @[Unit.scala 68:37]
  wire [15:0] BN_Array_8_io_input; // @[Unit.scala 68:37]
  wire [1:0] BN_Array_8_io_control; // @[Unit.scala 68:37]
  wire [15:0] BN_Array_8_io_output; // @[Unit.scala 68:37]
  wire  BN_Array_9_clock; // @[Unit.scala 68:37]
  wire  BN_Array_9_reset; // @[Unit.scala 68:37]
  wire [15:0] BN_Array_9_io_input; // @[Unit.scala 68:37]
  wire [1:0] BN_Array_9_io_control; // @[Unit.scala 68:37]
  wire [15:0] BN_Array_9_io_output; // @[Unit.scala 68:37]
  wire  BN_Array_10_clock; // @[Unit.scala 68:37]
  wire  BN_Array_10_reset; // @[Unit.scala 68:37]
  wire [15:0] BN_Array_10_io_input; // @[Unit.scala 68:37]
  wire [1:0] BN_Array_10_io_control; // @[Unit.scala 68:37]
  wire [15:0] BN_Array_10_io_output; // @[Unit.scala 68:37]
  wire  BN_Array_11_clock; // @[Unit.scala 68:37]
  wire  BN_Array_11_reset; // @[Unit.scala 68:37]
  wire [15:0] BN_Array_11_io_input; // @[Unit.scala 68:37]
  wire [1:0] BN_Array_11_io_control; // @[Unit.scala 68:37]
  wire [15:0] BN_Array_11_io_output; // @[Unit.scala 68:37]
  BN_Unit BN_Array_0 ( // @[Unit.scala 68:37]
    .clock(BN_Array_0_clock),
    .reset(BN_Array_0_reset),
    .io_input(BN_Array_0_io_input),
    .io_control(BN_Array_0_io_control),
    .io_output(BN_Array_0_io_output)
  );
  BN_Unit BN_Array_1 ( // @[Unit.scala 68:37]
    .clock(BN_Array_1_clock),
    .reset(BN_Array_1_reset),
    .io_input(BN_Array_1_io_input),
    .io_control(BN_Array_1_io_control),
    .io_output(BN_Array_1_io_output)
  );
  BN_Unit BN_Array_2 ( // @[Unit.scala 68:37]
    .clock(BN_Array_2_clock),
    .reset(BN_Array_2_reset),
    .io_input(BN_Array_2_io_input),
    .io_control(BN_Array_2_io_control),
    .io_output(BN_Array_2_io_output)
  );
  BN_Unit BN_Array_3 ( // @[Unit.scala 68:37]
    .clock(BN_Array_3_clock),
    .reset(BN_Array_3_reset),
    .io_input(BN_Array_3_io_input),
    .io_control(BN_Array_3_io_control),
    .io_output(BN_Array_3_io_output)
  );
  BN_Unit BN_Array_4 ( // @[Unit.scala 68:37]
    .clock(BN_Array_4_clock),
    .reset(BN_Array_4_reset),
    .io_input(BN_Array_4_io_input),
    .io_control(BN_Array_4_io_control),
    .io_output(BN_Array_4_io_output)
  );
  BN_Unit BN_Array_5 ( // @[Unit.scala 68:37]
    .clock(BN_Array_5_clock),
    .reset(BN_Array_5_reset),
    .io_input(BN_Array_5_io_input),
    .io_control(BN_Array_5_io_control),
    .io_output(BN_Array_5_io_output)
  );
  BN_Unit BN_Array_6 ( // @[Unit.scala 68:37]
    .clock(BN_Array_6_clock),
    .reset(BN_Array_6_reset),
    .io_input(BN_Array_6_io_input),
    .io_control(BN_Array_6_io_control),
    .io_output(BN_Array_6_io_output)
  );
  BN_Unit BN_Array_7 ( // @[Unit.scala 68:37]
    .clock(BN_Array_7_clock),
    .reset(BN_Array_7_reset),
    .io_input(BN_Array_7_io_input),
    .io_control(BN_Array_7_io_control),
    .io_output(BN_Array_7_io_output)
  );
  BN_Unit BN_Array_8 ( // @[Unit.scala 68:37]
    .clock(BN_Array_8_clock),
    .reset(BN_Array_8_reset),
    .io_input(BN_Array_8_io_input),
    .io_control(BN_Array_8_io_control),
    .io_output(BN_Array_8_io_output)
  );
  BN_Unit BN_Array_9 ( // @[Unit.scala 68:37]
    .clock(BN_Array_9_clock),
    .reset(BN_Array_9_reset),
    .io_input(BN_Array_9_io_input),
    .io_control(BN_Array_9_io_control),
    .io_output(BN_Array_9_io_output)
  );
  BN_Unit BN_Array_10 ( // @[Unit.scala 68:37]
    .clock(BN_Array_10_clock),
    .reset(BN_Array_10_reset),
    .io_input(BN_Array_10_io_input),
    .io_control(BN_Array_10_io_control),
    .io_output(BN_Array_10_io_output)
  );
  BN_Unit BN_Array_11 ( // @[Unit.scala 68:37]
    .clock(BN_Array_11_clock),
    .reset(BN_Array_11_reset),
    .io_input(BN_Array_11_io_input),
    .io_control(BN_Array_11_io_control),
    .io_output(BN_Array_11_io_output)
  );
  assign io_to_Relu6_0 = BN_Array_0_io_output; // @[Unit.scala 77:20]
  assign io_to_Relu6_1 = BN_Array_1_io_output; // @[Unit.scala 77:20]
  assign io_to_Relu6_2 = BN_Array_2_io_output; // @[Unit.scala 77:20]
  assign io_to_Relu6_3 = BN_Array_3_io_output; // @[Unit.scala 77:20]
  assign io_to_Relu6_4 = BN_Array_4_io_output; // @[Unit.scala 77:20]
  assign io_to_Relu6_5 = BN_Array_5_io_output; // @[Unit.scala 77:20]
  assign io_to_Relu6_6 = BN_Array_6_io_output; // @[Unit.scala 77:20]
  assign io_to_Relu6_7 = BN_Array_7_io_output; // @[Unit.scala 77:20]
  assign io_to_Relu6_8 = BN_Array_8_io_output; // @[Unit.scala 77:20]
  assign io_to_Relu6_9 = BN_Array_9_io_output; // @[Unit.scala 77:20]
  assign io_to_Relu6_10 = BN_Array_10_io_output; // @[Unit.scala 77:20]
  assign io_to_Relu6_11 = BN_Array_11_io_output; // @[Unit.scala 77:20]
  assign BN_Array_0_clock = clock;
  assign BN_Array_0_reset = reset;
  assign BN_Array_0_io_input = io_from_PE_0; // @[Unit.scala 72:26]
  assign BN_Array_0_io_control = io_control_0; // @[Unit.scala 73:28]
  assign BN_Array_1_clock = clock;
  assign BN_Array_1_reset = reset;
  assign BN_Array_1_io_input = io_from_PE_1; // @[Unit.scala 72:26]
  assign BN_Array_1_io_control = io_control_1; // @[Unit.scala 73:28]
  assign BN_Array_2_clock = clock;
  assign BN_Array_2_reset = reset;
  assign BN_Array_2_io_input = io_from_PE_2; // @[Unit.scala 72:26]
  assign BN_Array_2_io_control = io_control_2; // @[Unit.scala 73:28]
  assign BN_Array_3_clock = clock;
  assign BN_Array_3_reset = reset;
  assign BN_Array_3_io_input = io_from_PE_3; // @[Unit.scala 72:26]
  assign BN_Array_3_io_control = io_control_3; // @[Unit.scala 73:28]
  assign BN_Array_4_clock = clock;
  assign BN_Array_4_reset = reset;
  assign BN_Array_4_io_input = io_from_PE_4; // @[Unit.scala 72:26]
  assign BN_Array_4_io_control = io_control_4; // @[Unit.scala 73:28]
  assign BN_Array_5_clock = clock;
  assign BN_Array_5_reset = reset;
  assign BN_Array_5_io_input = io_from_PE_5; // @[Unit.scala 72:26]
  assign BN_Array_5_io_control = io_control_5; // @[Unit.scala 73:28]
  assign BN_Array_6_clock = clock;
  assign BN_Array_6_reset = reset;
  assign BN_Array_6_io_input = io_from_PE_6; // @[Unit.scala 72:26]
  assign BN_Array_6_io_control = io_control_6; // @[Unit.scala 73:28]
  assign BN_Array_7_clock = clock;
  assign BN_Array_7_reset = reset;
  assign BN_Array_7_io_input = io_from_PE_7; // @[Unit.scala 72:26]
  assign BN_Array_7_io_control = io_control_7; // @[Unit.scala 73:28]
  assign BN_Array_8_clock = clock;
  assign BN_Array_8_reset = reset;
  assign BN_Array_8_io_input = io_from_PE_8; // @[Unit.scala 72:26]
  assign BN_Array_8_io_control = io_control_8; // @[Unit.scala 73:28]
  assign BN_Array_9_clock = clock;
  assign BN_Array_9_reset = reset;
  assign BN_Array_9_io_input = io_from_PE_9; // @[Unit.scala 72:26]
  assign BN_Array_9_io_control = io_control_9; // @[Unit.scala 73:28]
  assign BN_Array_10_clock = clock;
  assign BN_Array_10_reset = reset;
  assign BN_Array_10_io_input = io_from_PE_10; // @[Unit.scala 72:26]
  assign BN_Array_10_io_control = io_control_10; // @[Unit.scala 73:28]
  assign BN_Array_11_clock = clock;
  assign BN_Array_11_reset = reset;
  assign BN_Array_11_io_input = io_from_PE_11; // @[Unit.scala 72:26]
  assign BN_Array_11_io_control = io_control_11; // @[Unit.scala 73:28]
endmodule
module Relu6_Unit(
  input  [15:0] io_input,
  input         io_control,
  output [15:0] io_output
);
  wire [15:0] _GEN_0 = ~io_input[15] & io_input <= 16'h4600 ? io_input : 16'h4600; // @[Unit.scala 97:72 Unit.scala 98:17 Unit.scala 101:17]
  wire [15:0] _GEN_1 = io_input[15] ? 16'h0 : _GEN_0; // @[Unit.scala 94:38 Unit.scala 95:17]
  assign io_output = ~io_control ? io_input : _GEN_1; // @[Unit.scala 89:27 Unit.scala 90:15]
endmodule
module Relu6_Unit_Array(
  input  [15:0] io_input_0,
  input  [15:0] io_input_1,
  input  [15:0] io_input_2,
  input  [15:0] io_input_3,
  input  [15:0] io_input_4,
  input  [15:0] io_input_5,
  input  [15:0] io_input_6,
  input  [15:0] io_input_7,
  input  [15:0] io_input_8,
  input  [15:0] io_input_9,
  input  [15:0] io_input_10,
  input  [15:0] io_input_11,
  input         io_control_0,
  input         io_control_1,
  input         io_control_2,
  input         io_control_3,
  input         io_control_4,
  input         io_control_5,
  input         io_control_6,
  input         io_control_7,
  input         io_control_8,
  input         io_control_9,
  input         io_control_10,
  input         io_control_11,
  output [15:0] io_output_0,
  output [15:0] io_output_1,
  output [15:0] io_output_2,
  output [15:0] io_output_3,
  output [15:0] io_output_4,
  output [15:0] io_output_5,
  output [15:0] io_output_6,
  output [15:0] io_output_7,
  output [15:0] io_output_8,
  output [15:0] io_output_9,
  output [15:0] io_output_10,
  output [15:0] io_output_11
);
  wire [15:0] Relu6_Array_0_io_input; // @[Unit.scala 114:40]
  wire  Relu6_Array_0_io_control; // @[Unit.scala 114:40]
  wire [15:0] Relu6_Array_0_io_output; // @[Unit.scala 114:40]
  wire [15:0] Relu6_Array_1_io_input; // @[Unit.scala 114:40]
  wire  Relu6_Array_1_io_control; // @[Unit.scala 114:40]
  wire [15:0] Relu6_Array_1_io_output; // @[Unit.scala 114:40]
  wire [15:0] Relu6_Array_2_io_input; // @[Unit.scala 114:40]
  wire  Relu6_Array_2_io_control; // @[Unit.scala 114:40]
  wire [15:0] Relu6_Array_2_io_output; // @[Unit.scala 114:40]
  wire [15:0] Relu6_Array_3_io_input; // @[Unit.scala 114:40]
  wire  Relu6_Array_3_io_control; // @[Unit.scala 114:40]
  wire [15:0] Relu6_Array_3_io_output; // @[Unit.scala 114:40]
  wire [15:0] Relu6_Array_4_io_input; // @[Unit.scala 114:40]
  wire  Relu6_Array_4_io_control; // @[Unit.scala 114:40]
  wire [15:0] Relu6_Array_4_io_output; // @[Unit.scala 114:40]
  wire [15:0] Relu6_Array_5_io_input; // @[Unit.scala 114:40]
  wire  Relu6_Array_5_io_control; // @[Unit.scala 114:40]
  wire [15:0] Relu6_Array_5_io_output; // @[Unit.scala 114:40]
  wire [15:0] Relu6_Array_6_io_input; // @[Unit.scala 114:40]
  wire  Relu6_Array_6_io_control; // @[Unit.scala 114:40]
  wire [15:0] Relu6_Array_6_io_output; // @[Unit.scala 114:40]
  wire [15:0] Relu6_Array_7_io_input; // @[Unit.scala 114:40]
  wire  Relu6_Array_7_io_control; // @[Unit.scala 114:40]
  wire [15:0] Relu6_Array_7_io_output; // @[Unit.scala 114:40]
  wire [15:0] Relu6_Array_8_io_input; // @[Unit.scala 114:40]
  wire  Relu6_Array_8_io_control; // @[Unit.scala 114:40]
  wire [15:0] Relu6_Array_8_io_output; // @[Unit.scala 114:40]
  wire [15:0] Relu6_Array_9_io_input; // @[Unit.scala 114:40]
  wire  Relu6_Array_9_io_control; // @[Unit.scala 114:40]
  wire [15:0] Relu6_Array_9_io_output; // @[Unit.scala 114:40]
  wire [15:0] Relu6_Array_10_io_input; // @[Unit.scala 114:40]
  wire  Relu6_Array_10_io_control; // @[Unit.scala 114:40]
  wire [15:0] Relu6_Array_10_io_output; // @[Unit.scala 114:40]
  wire [15:0] Relu6_Array_11_io_input; // @[Unit.scala 114:40]
  wire  Relu6_Array_11_io_control; // @[Unit.scala 114:40]
  wire [15:0] Relu6_Array_11_io_output; // @[Unit.scala 114:40]
  Relu6_Unit Relu6_Array_0 ( // @[Unit.scala 114:40]
    .io_input(Relu6_Array_0_io_input),
    .io_control(Relu6_Array_0_io_control),
    .io_output(Relu6_Array_0_io_output)
  );
  Relu6_Unit Relu6_Array_1 ( // @[Unit.scala 114:40]
    .io_input(Relu6_Array_1_io_input),
    .io_control(Relu6_Array_1_io_control),
    .io_output(Relu6_Array_1_io_output)
  );
  Relu6_Unit Relu6_Array_2 ( // @[Unit.scala 114:40]
    .io_input(Relu6_Array_2_io_input),
    .io_control(Relu6_Array_2_io_control),
    .io_output(Relu6_Array_2_io_output)
  );
  Relu6_Unit Relu6_Array_3 ( // @[Unit.scala 114:40]
    .io_input(Relu6_Array_3_io_input),
    .io_control(Relu6_Array_3_io_control),
    .io_output(Relu6_Array_3_io_output)
  );
  Relu6_Unit Relu6_Array_4 ( // @[Unit.scala 114:40]
    .io_input(Relu6_Array_4_io_input),
    .io_control(Relu6_Array_4_io_control),
    .io_output(Relu6_Array_4_io_output)
  );
  Relu6_Unit Relu6_Array_5 ( // @[Unit.scala 114:40]
    .io_input(Relu6_Array_5_io_input),
    .io_control(Relu6_Array_5_io_control),
    .io_output(Relu6_Array_5_io_output)
  );
  Relu6_Unit Relu6_Array_6 ( // @[Unit.scala 114:40]
    .io_input(Relu6_Array_6_io_input),
    .io_control(Relu6_Array_6_io_control),
    .io_output(Relu6_Array_6_io_output)
  );
  Relu6_Unit Relu6_Array_7 ( // @[Unit.scala 114:40]
    .io_input(Relu6_Array_7_io_input),
    .io_control(Relu6_Array_7_io_control),
    .io_output(Relu6_Array_7_io_output)
  );
  Relu6_Unit Relu6_Array_8 ( // @[Unit.scala 114:40]
    .io_input(Relu6_Array_8_io_input),
    .io_control(Relu6_Array_8_io_control),
    .io_output(Relu6_Array_8_io_output)
  );
  Relu6_Unit Relu6_Array_9 ( // @[Unit.scala 114:40]
    .io_input(Relu6_Array_9_io_input),
    .io_control(Relu6_Array_9_io_control),
    .io_output(Relu6_Array_9_io_output)
  );
  Relu6_Unit Relu6_Array_10 ( // @[Unit.scala 114:40]
    .io_input(Relu6_Array_10_io_input),
    .io_control(Relu6_Array_10_io_control),
    .io_output(Relu6_Array_10_io_output)
  );
  Relu6_Unit Relu6_Array_11 ( // @[Unit.scala 114:40]
    .io_input(Relu6_Array_11_io_input),
    .io_control(Relu6_Array_11_io_control),
    .io_output(Relu6_Array_11_io_output)
  );
  assign io_output_0 = Relu6_Array_0_io_output; // @[Unit.scala 120:18]
  assign io_output_1 = Relu6_Array_1_io_output; // @[Unit.scala 120:18]
  assign io_output_2 = Relu6_Array_2_io_output; // @[Unit.scala 120:18]
  assign io_output_3 = Relu6_Array_3_io_output; // @[Unit.scala 120:18]
  assign io_output_4 = Relu6_Array_4_io_output; // @[Unit.scala 120:18]
  assign io_output_5 = Relu6_Array_5_io_output; // @[Unit.scala 120:18]
  assign io_output_6 = Relu6_Array_6_io_output; // @[Unit.scala 120:18]
  assign io_output_7 = Relu6_Array_7_io_output; // @[Unit.scala 120:18]
  assign io_output_8 = Relu6_Array_8_io_output; // @[Unit.scala 120:18]
  assign io_output_9 = Relu6_Array_9_io_output; // @[Unit.scala 120:18]
  assign io_output_10 = Relu6_Array_10_io_output; // @[Unit.scala 120:18]
  assign io_output_11 = Relu6_Array_11_io_output; // @[Unit.scala 120:18]
  assign Relu6_Array_0_io_input = io_input_0; // @[Unit.scala 118:29]
  assign Relu6_Array_0_io_control = io_control_0; // @[Unit.scala 119:31]
  assign Relu6_Array_1_io_input = io_input_1; // @[Unit.scala 118:29]
  assign Relu6_Array_1_io_control = io_control_1; // @[Unit.scala 119:31]
  assign Relu6_Array_2_io_input = io_input_2; // @[Unit.scala 118:29]
  assign Relu6_Array_2_io_control = io_control_2; // @[Unit.scala 119:31]
  assign Relu6_Array_3_io_input = io_input_3; // @[Unit.scala 118:29]
  assign Relu6_Array_3_io_control = io_control_3; // @[Unit.scala 119:31]
  assign Relu6_Array_4_io_input = io_input_4; // @[Unit.scala 118:29]
  assign Relu6_Array_4_io_control = io_control_4; // @[Unit.scala 119:31]
  assign Relu6_Array_5_io_input = io_input_5; // @[Unit.scala 118:29]
  assign Relu6_Array_5_io_control = io_control_5; // @[Unit.scala 119:31]
  assign Relu6_Array_6_io_input = io_input_6; // @[Unit.scala 118:29]
  assign Relu6_Array_6_io_control = io_control_6; // @[Unit.scala 119:31]
  assign Relu6_Array_7_io_input = io_input_7; // @[Unit.scala 118:29]
  assign Relu6_Array_7_io_control = io_control_7; // @[Unit.scala 119:31]
  assign Relu6_Array_8_io_input = io_input_8; // @[Unit.scala 118:29]
  assign Relu6_Array_8_io_control = io_control_8; // @[Unit.scala 119:31]
  assign Relu6_Array_9_io_input = io_input_9; // @[Unit.scala 118:29]
  assign Relu6_Array_9_io_control = io_control_9; // @[Unit.scala 119:31]
  assign Relu6_Array_10_io_input = io_input_10; // @[Unit.scala 118:29]
  assign Relu6_Array_10_io_control = io_control_10; // @[Unit.scala 119:31]
  assign Relu6_Array_11_io_input = io_input_11; // @[Unit.scala 118:29]
  assign Relu6_Array_11_io_control = io_control_11; // @[Unit.scala 119:31]
endmodule
module activation_Unit(
  input         clock,
  input         reset,
  input  [15:0] io_input,
  input  [1:0]  io_control,
  output [15:0] io_output
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] relu6_io_input; // @[Unit.scala 132:21]
  wire  relu6_io_control; // @[Unit.scala 132:21]
  wire [15:0] relu6_io_output; // @[Unit.scala 132:21]
  wire [15:0] FP16MAC_io_a; // @[Unit.scala 137:23]
  wire [15:0] FP16MAC_io_b; // @[Unit.scala 137:23]
  wire [15:0] FP16MAC_io_c; // @[Unit.scala 137:23]
  wire [15:0] FP16MAC_io_out; // @[Unit.scala 137:23]
  reg [15:0] output_reg; // @[Unit.scala 143:27]
  wire  _T_53 = ~io_input[15]; // @[Unit.scala 208:36]
  wire [15:0] _GEN_0 = _T_53 & io_input > 16'h4700 & io_input <= 16'h4800 ? io_input : 16'h0; // @[Unit.scala 250:99 Unit.scala 251:20 Unit.scala 257:22]
  wire [12:0] _GEN_1 = _T_53 & io_input > 16'h4700 & io_input <= 16'h4800 ? 13'h10ea : 13'h0; // @[Unit.scala 250:99 Unit.scala 252:20 Unit.scala 258:22]
  wire [13:0] _GEN_2 = _T_53 & io_input > 16'h4700 & io_input <= 16'h4800 ? 14'h3bf6 : 14'h0; // @[Unit.scala 250:99 Unit.scala 253:20 Unit.scala 259:22]
  wire [15:0] _GEN_3 = _T_53 & io_input > 16'h4700 & io_input <= 16'h4800 ? FP16MAC_io_out : 16'h3c00; // @[Unit.scala 250:99 Unit.scala 254:18 Unit.scala 260:20]
  wire [15:0] _GEN_4 = _T_53 & io_input > 16'h4600 & io_input <= 16'h4700 ? io_input : _GEN_0; // @[Unit.scala 244:98 Unit.scala 245:20]
  wire [12:0] _GEN_5 = _T_53 & io_input > 16'h4600 & io_input <= 16'h4700 ? 13'h1624 : _GEN_1; // @[Unit.scala 244:98 Unit.scala 246:20]
  wire [13:0] _GEN_6 = _T_53 & io_input > 16'h4600 & io_input <= 16'h4700 ? 14'h3be8 : _GEN_2; // @[Unit.scala 244:98 Unit.scala 247:20]
  wire [15:0] _GEN_7 = _T_53 & io_input > 16'h4600 & io_input <= 16'h4700 ? FP16MAC_io_out : _GEN_3; // @[Unit.scala 244:98 Unit.scala 248:18]
  wire [15:0] _GEN_8 = _T_53 & io_input > 16'h4500 & io_input <= 16'h4600 ? io_input : _GEN_4; // @[Unit.scala 238:98 Unit.scala 239:20]
  wire [12:0] _GEN_9 = _T_53 & io_input > 16'h4500 & io_input <= 16'h4600 ? 13'h1c4d : _GEN_5; // @[Unit.scala 238:98 Unit.scala 240:20]
  wire [13:0] _GEN_10 = _T_53 & io_input > 16'h4500 & io_input <= 16'h4600 ? 14'h3bc8 : _GEN_6; // @[Unit.scala 238:98 Unit.scala 241:20]
  wire [15:0] _GEN_11 = _T_53 & io_input > 16'h4500 & io_input <= 16'h4600 ? FP16MAC_io_out : _GEN_7; // @[Unit.scala 238:98 Unit.scala 242:18]
  wire [15:0] _GEN_12 = _T_53 & io_input > 16'h4400 & io_input <= 16'h4500 ? io_input : _GEN_8; // @[Unit.scala 232:98 Unit.scala 233:20]
  wire [13:0] _GEN_13 = _T_53 & io_input > 16'h4400 & io_input <= 16'h4500 ? 14'h21ae : {{1'd0}, _GEN_9}; // @[Unit.scala 232:98 Unit.scala 234:20]
  wire [13:0] _GEN_14 = _T_53 & io_input > 16'h4400 & io_input <= 16'h4500 ? 14'h3b82 : _GEN_10; // @[Unit.scala 232:98 Unit.scala 235:20]
  wire [15:0] _GEN_15 = _T_53 & io_input > 16'h4400 & io_input <= 16'h4500 ? FP16MAC_io_out : _GEN_11; // @[Unit.scala 232:98 Unit.scala 236:18]
  wire [15:0] _GEN_16 = _T_53 & io_input > 16'h4200 & io_input <= 16'h4400 ? io_input : _GEN_12; // @[Unit.scala 226:98 Unit.scala 227:20]
  wire [13:0] _GEN_17 = _T_53 & io_input > 16'h4200 & io_input <= 16'h4400 ? 14'h2773 : _GEN_13; // @[Unit.scala 226:98 Unit.scala 228:20]
  wire [13:0] _GEN_18 = _T_53 & io_input > 16'h4200 & io_input <= 16'h4400 ? 14'h3af1 : _GEN_14; // @[Unit.scala 226:98 Unit.scala 229:20]
  wire [15:0] _GEN_19 = _T_53 & io_input > 16'h4200 & io_input <= 16'h4400 ? FP16MAC_io_out : _GEN_15; // @[Unit.scala 226:98 Unit.scala 230:18]
  wire [15:0] _GEN_20 = _T_53 & io_input > 16'h4000 & io_input <= 16'h4200 ? io_input : _GEN_16; // @[Unit.scala 220:98 Unit.scala 221:20]
  wire [13:0] _GEN_21 = _T_53 & io_input > 16'h4000 & io_input <= 16'h4200 ? 14'h2c8c : _GEN_17; // @[Unit.scala 220:98 Unit.scala 222:20]
  wire [13:0] _GEN_22 = _T_53 & io_input > 16'h4000 & io_input <= 16'h4200 ? 14'h39f3 : _GEN_18; // @[Unit.scala 220:98 Unit.scala 223:20]
  wire [15:0] _GEN_23 = _T_53 & io_input > 16'h4000 & io_input <= 16'h4200 ? FP16MAC_io_out : _GEN_19; // @[Unit.scala 220:98 Unit.scala 224:18]
  wire [15:0] _GEN_24 = _T_53 & io_input > 16'h3c00 & io_input <= 16'h4000 ? io_input : _GEN_20; // @[Unit.scala 214:98 Unit.scala 215:20]
  wire [13:0] _GEN_25 = _T_53 & io_input > 16'h3c00 & io_input <= 16'h4000 ? 14'h30c8 : _GEN_21; // @[Unit.scala 214:98 Unit.scala 216:20]
  wire [13:0] _GEN_26 = _T_53 & io_input > 16'h3c00 & io_input <= 16'h4000 ? 14'h38b6 : _GEN_22; // @[Unit.scala 214:98 Unit.scala 217:20]
  wire [15:0] _GEN_27 = _T_53 & io_input > 16'h3c00 & io_input <= 16'h4000 ? FP16MAC_io_out : _GEN_23; // @[Unit.scala 214:98 Unit.scala 218:18]
  wire [15:0] _GEN_28 = ~io_input[15] & io_input <= 16'h3c00 ? io_input : _GEN_24; // @[Unit.scala 208:93 Unit.scala 209:20]
  wire [13:0] _GEN_29 = ~io_input[15] & io_input <= 16'h3c00 ? 14'h3371 : _GEN_25; // @[Unit.scala 208:93 Unit.scala 210:20]
  wire [13:0] _GEN_30 = ~io_input[15] & io_input <= 16'h3c00 ? 14'h3807 : _GEN_26; // @[Unit.scala 208:93 Unit.scala 211:20]
  wire [15:0] _GEN_31 = ~io_input[15] & io_input <= 16'h3c00 ? FP16MAC_io_out : _GEN_27; // @[Unit.scala 208:93 Unit.scala 212:18]
  wire [15:0] _GEN_32 = io_input[15] & io_input < 16'hbc00 ? io_input : _GEN_28; // @[Unit.scala 202:71 Unit.scala 203:20]
  wire [13:0] _GEN_33 = io_input[15] & io_input < 16'hbc00 ? 14'h3371 : _GEN_29; // @[Unit.scala 202:71 Unit.scala 204:20]
  wire [13:0] _GEN_34 = io_input[15] & io_input < 16'hbc00 ? 14'h37f0 : _GEN_30; // @[Unit.scala 202:71 Unit.scala 205:20]
  wire [15:0] _GEN_35 = io_input[15] & io_input < 16'hbc00 ? FP16MAC_io_out : _GEN_31; // @[Unit.scala 202:71 Unit.scala 206:18]
  wire [15:0] _GEN_36 = io_input[15] & io_input < 16'hc000 & io_input >= 16'hbc00 ? io_input : _GEN_32; // @[Unit.scala 196:98 Unit.scala 197:20]
  wire [13:0] _GEN_37 = io_input[15] & io_input < 16'hc000 & io_input >= 16'hbc00 ? 14'h30c8 : _GEN_33; // @[Unit.scala 196:98 Unit.scala 198:20]
  wire [13:0] _GEN_38 = io_input[15] & io_input < 16'hc000 & io_input >= 16'hbc00 ? 14'h3692 : _GEN_34; // @[Unit.scala 196:98 Unit.scala 199:20]
  wire [15:0] _GEN_39 = io_input[15] & io_input < 16'hc000 & io_input >= 16'hbc00 ? FP16MAC_io_out : _GEN_35; // @[Unit.scala 196:98 Unit.scala 200:18]
  wire [15:0] _GEN_40 = io_input[15] & io_input < 16'hc200 & io_input >= 16'hc000 ? io_input : _GEN_36; // @[Unit.scala 190:98 Unit.scala 191:20]
  wire [13:0] _GEN_41 = io_input[15] & io_input < 16'hc200 & io_input >= 16'hc000 ? 14'h2c8c : _GEN_37; // @[Unit.scala 190:98 Unit.scala 192:20]
  wire [13:0] _GEN_42 = io_input[15] & io_input < 16'hc200 & io_input >= 16'hc000 ? 14'h3419 : _GEN_38; // @[Unit.scala 190:98 Unit.scala 193:20]
  wire [15:0] _GEN_43 = io_input[15] & io_input < 16'hc200 & io_input >= 16'hc000 ? FP16MAC_io_out : _GEN_39; // @[Unit.scala 190:98 Unit.scala 194:18]
  wire [15:0] _GEN_44 = io_input[15] & io_input < 16'hc400 & io_input >= 16'hc200 ? io_input : _GEN_40; // @[Unit.scala 184:98 Unit.scala 185:20]
  wire [13:0] _GEN_45 = io_input[15] & io_input < 16'hc400 & io_input >= 16'hc200 ? 14'h2773 : _GEN_41; // @[Unit.scala 184:98 Unit.scala 186:20]
  wire [13:0] _GEN_46 = io_input[15] & io_input < 16'hc400 & io_input >= 16'hc200 ? 14'h303a : _GEN_42; // @[Unit.scala 184:98 Unit.scala 187:20]
  wire [15:0] _GEN_47 = io_input[15] & io_input < 16'hc400 & io_input >= 16'hc200 ? FP16MAC_io_out : _GEN_43; // @[Unit.scala 184:98 Unit.scala 188:18]
  wire [15:0] _GEN_48 = io_input[15] & io_input < 16'hc500 & io_input >= 16'hc400 ? io_input : _GEN_44; // @[Unit.scala 178:98 Unit.scala 179:20]
  wire [13:0] _GEN_49 = io_input[15] & io_input < 16'hc500 & io_input >= 16'hc400 ? 14'h21ae : _GEN_45; // @[Unit.scala 178:98 Unit.scala 180:20]
  wire [13:0] _GEN_50 = io_input[15] & io_input < 16'hc500 & io_input >= 16'hc400 ? 14'h2bdf : _GEN_46; // @[Unit.scala 178:98 Unit.scala 181:20]
  wire [15:0] _GEN_51 = io_input[15] & io_input < 16'hc500 & io_input >= 16'hc400 ? FP16MAC_io_out : _GEN_47; // @[Unit.scala 178:98 Unit.scala 182:18]
  wire [15:0] _GEN_52 = io_input[15] & io_input < 16'hc600 & io_input >= 16'hc500 ? io_input : _GEN_48; // @[Unit.scala 172:98 Unit.scala 173:20]
  wire [13:0] _GEN_53 = io_input[15] & io_input < 16'hc600 & io_input >= 16'hc500 ? 14'h1c4d : _GEN_49; // @[Unit.scala 172:98 Unit.scala 174:20]
  wire [13:0] _GEN_54 = io_input[15] & io_input < 16'hc600 & io_input >= 16'hc500 ? 14'h26f0 : _GEN_50; // @[Unit.scala 172:98 Unit.scala 175:20]
  wire [15:0] _GEN_55 = io_input[15] & io_input < 16'hc600 & io_input >= 16'hc500 ? FP16MAC_io_out : _GEN_51; // @[Unit.scala 172:98 Unit.scala 176:18]
  wire [15:0] _GEN_56 = io_input[15] & io_input < 16'hc700 & io_input >= 16'hc600 ? io_input : _GEN_52; // @[Unit.scala 166:98 Unit.scala 167:20]
  wire [13:0] _GEN_57 = io_input[15] & io_input < 16'hc700 & io_input >= 16'hc600 ? 14'h1624 : _GEN_53; // @[Unit.scala 166:98 Unit.scala 168:20]
  wire [13:0] _GEN_58 = io_input[15] & io_input < 16'hc700 & io_input >= 16'hc600 ? 14'h21f0 : _GEN_54; // @[Unit.scala 166:98 Unit.scala 169:20]
  wire [15:0] _GEN_59 = io_input[15] & io_input < 16'hc700 & io_input >= 16'hc600 ? FP16MAC_io_out : _GEN_55; // @[Unit.scala 166:98 Unit.scala 170:18]
  wire [15:0] _GEN_60 = io_input[15] & io_input < 16'hc800 & io_input >= 16'hc700 ? io_input : _GEN_56; // @[Unit.scala 160:98 Unit.scala 161:20]
  wire [13:0] _GEN_61 = io_input[15] & io_input < 16'hc800 & io_input >= 16'hc700 ? 14'h1e24 : _GEN_57; // @[Unit.scala 160:98 Unit.scala 162:20]
  wire [13:0] _GEN_62 = io_input[15] & io_input < 16'hc800 & io_input >= 16'hc700 ? 14'h1cea : _GEN_58; // @[Unit.scala 160:98 Unit.scala 163:20]
  wire [15:0] _GEN_63 = io_input[15] & io_input < 16'hc800 & io_input >= 16'hc700 ? FP16MAC_io_out : _GEN_59; // @[Unit.scala 160:98 Unit.scala 164:18]
  wire [15:0] _GEN_64 = io_input[15] & io_input >= 16'hc800 ? 16'h0 : _GEN_60; // @[Unit.scala 154:67 Unit.scala 155:20]
  wire [13:0] _GEN_65 = io_input[15] & io_input >= 16'hc800 ? 14'h0 : _GEN_61; // @[Unit.scala 154:67 Unit.scala 156:20]
  wire [13:0] _GEN_66 = io_input[15] & io_input >= 16'hc800 ? 14'h0 : _GEN_62; // @[Unit.scala 154:67 Unit.scala 157:20]
  wire [15:0] _GEN_70 = io_control == 2'h1 ? _GEN_64 : 16'h0; // @[Unit.scala 153:32]
  wire [13:0] _GEN_71 = io_control == 2'h1 ? _GEN_65 : 14'h0; // @[Unit.scala 153:32]
  wire [13:0] _GEN_72 = io_control == 2'h1 ? _GEN_66 : 14'h0; // @[Unit.scala 153:32]
  wire [13:0] _GEN_75 = io_control == 2'h0 ? 14'h0 : _GEN_71; // @[Unit.scala 146:27 Unit.scala 148:18]
  wire [13:0] _GEN_76 = io_control == 2'h0 ? 14'h0 : _GEN_72; // @[Unit.scala 146:27 Unit.scala 149:18]
  Relu6_Unit relu6 ( // @[Unit.scala 132:21]
    .io_input(relu6_io_input),
    .io_control(relu6_io_control),
    .io_output(relu6_io_output)
  );
  FP16MulAdder FP16MAC ( // @[Unit.scala 137:23]
    .io_a(FP16MAC_io_a),
    .io_b(FP16MAC_io_b),
    .io_c(FP16MAC_io_c),
    .io_out(FP16MAC_io_out)
  );
  assign io_output = output_reg; // @[Unit.scala 144:13]
  assign relu6_io_input = io_input; // @[Unit.scala 134:18]
  assign relu6_io_control = 1'h1; // @[Unit.scala 133:20]
  assign FP16MAC_io_a = io_control == 2'h0 ? 16'h0 : _GEN_70; // @[Unit.scala 146:27 Unit.scala 147:18]
  assign FP16MAC_io_b = {{2'd0}, _GEN_75}; // @[Unit.scala 146:27 Unit.scala 148:18]
  assign FP16MAC_io_c = {{2'd0}, _GEN_76}; // @[Unit.scala 146:27 Unit.scala 149:18]
  always @(posedge clock) begin
    if (reset) begin // @[Unit.scala 143:27]
      output_reg <= 16'h0; // @[Unit.scala 143:27]
    end else if (io_control == 2'h0) begin // @[Unit.scala 146:27]
      output_reg <= io_input; // @[Unit.scala 150:16]
    end else if (io_control == 2'h1) begin // @[Unit.scala 153:32]
      if (io_input[15] & io_input >= 16'hc800) begin // @[Unit.scala 154:67]
        output_reg <= 16'h0; // @[Unit.scala 158:18]
      end else begin
        output_reg <= _GEN_63;
      end
    end else if (io_control == 2'h2) begin // @[Unit.scala 264:32]
      output_reg <= io_input; // @[Unit.scala 265:16]
    end else begin
      output_reg <= relu6_io_output; // @[Unit.scala 272:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  output_reg = _RAND_0[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module accumulator_registers(
  input         clock,
  input         reset,
  input  [5:0]  io_rdAddr,
  output [15:0] io_rdData,
  input         io_wrEna,
  input  [15:0] io_wrData,
  input  [5:0]  io_wrAddr
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] FP16MAC_io_a; // @[Unit.scala 389:23]
  wire [15:0] FP16MAC_io_b; // @[Unit.scala 389:23]
  wire [15:0] FP16MAC_io_c; // @[Unit.scala 389:23]
  wire [15:0] FP16MAC_io_out; // @[Unit.scala 389:23]
  reg [15:0] register_0; // @[Unit.scala 386:25]
  reg [15:0] register_1; // @[Unit.scala 386:25]
  reg [15:0] register_2; // @[Unit.scala 386:25]
  reg [15:0] register_3; // @[Unit.scala 386:25]
  wire [15:0] _GEN_1 = 2'h1 == io_rdAddr[1:0] ? register_1 : register_0; // @[Unit.scala 394:13 Unit.scala 394:13]
  wire [15:0] _GEN_2 = 2'h2 == io_rdAddr[1:0] ? register_2 : _GEN_1; // @[Unit.scala 394:13 Unit.scala 394:13]
  wire [15:0] _GEN_5 = 2'h1 == io_wrAddr[1:0] ? register_1 : register_0; // @[Unit.scala 398:18 Unit.scala 398:18]
  wire [15:0] _GEN_6 = 2'h2 == io_wrAddr[1:0] ? register_2 : _GEN_5; // @[Unit.scala 398:18 Unit.scala 398:18]
  wire [15:0] _GEN_7 = 2'h3 == io_wrAddr[1:0] ? register_3 : _GEN_6; // @[Unit.scala 398:18 Unit.scala 398:18]
  wire [15:0] _register_T = FP16MAC_io_out; // @[Unit.scala 399:25 Unit.scala 399:25]
  wire [13:0] _GEN_13 = io_wrEna ? 14'h3c00 : 14'h0; // @[Unit.scala 395:17 Unit.scala 397:18 Unit.scala 403:20]
  FP16MulAdder FP16MAC ( // @[Unit.scala 389:23]
    .io_a(FP16MAC_io_a),
    .io_b(FP16MAC_io_b),
    .io_c(FP16MAC_io_c),
    .io_out(FP16MAC_io_out)
  );
  assign io_rdData = 2'h3 == io_rdAddr[1:0] ? register_3 : _GEN_2; // @[Unit.scala 394:13 Unit.scala 394:13]
  assign FP16MAC_io_a = io_wrEna ? io_wrData : 16'h0; // @[Unit.scala 395:17 Unit.scala 396:18 Unit.scala 402:20]
  assign FP16MAC_io_b = {{2'd0}, _GEN_13}; // @[Unit.scala 395:17 Unit.scala 397:18 Unit.scala 403:20]
  assign FP16MAC_io_c = io_wrEna ? _GEN_7 : 16'h0; // @[Unit.scala 395:17 Unit.scala 398:18 Unit.scala 404:20]
  always @(posedge clock) begin
    if (reset) begin // @[Unit.scala 386:25]
      register_0 <= 16'h0; // @[Unit.scala 386:25]
    end else if (io_wrEna) begin // @[Unit.scala 395:17]
      if (2'h0 == io_wrAddr[1:0]) begin // @[Unit.scala 399:25]
        register_0 <= _register_T; // @[Unit.scala 399:25]
      end
    end
    if (reset) begin // @[Unit.scala 386:25]
      register_1 <= 16'h0; // @[Unit.scala 386:25]
    end else if (io_wrEna) begin // @[Unit.scala 395:17]
      if (2'h1 == io_wrAddr[1:0]) begin // @[Unit.scala 399:25]
        register_1 <= _register_T; // @[Unit.scala 399:25]
      end
    end
    if (reset) begin // @[Unit.scala 386:25]
      register_2 <= 16'h0; // @[Unit.scala 386:25]
    end else if (io_wrEna) begin // @[Unit.scala 395:17]
      if (2'h2 == io_wrAddr[1:0]) begin // @[Unit.scala 399:25]
        register_2 <= _register_T; // @[Unit.scala 399:25]
      end
    end
    if (reset) begin // @[Unit.scala 386:25]
      register_3 <= 16'h0; // @[Unit.scala 386:25]
    end else if (io_wrEna) begin // @[Unit.scala 395:17]
      if (2'h3 == io_wrAddr[1:0]) begin // @[Unit.scala 399:25]
        register_3 <= _register_T; // @[Unit.scala 399:25]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  register_0 = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  register_1 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  register_2 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  register_3 = _RAND_3[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ht(
  input         clock,
  input         reset,
  output [15:0] io_to_PE_0,
  output [15:0] io_to_PE_1,
  output [15:0] io_to_PE_2,
  output [15:0] io_to_PE_3,
  output [15:0] io_to_PE_4,
  output [15:0] io_to_PE_5,
  output [15:0] io_to_PE_6,
  output [15:0] io_to_PE_7,
  output [15:0] io_to_PE_8,
  output [15:0] io_to_PE_9,
  output [15:0] io_to_PE_10,
  output [15:0] io_to_PE_11,
  input  [2:0]  io_to_PE_control,
  output [15:0] io_rdData,
  input         io_wrEna,
  input  [15:0] io_wrData,
  input  [5:0]  io_wrAddr
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] FP16MAC_io_a; // @[Unit.scala 422:23]
  wire [15:0] FP16MAC_io_b; // @[Unit.scala 422:23]
  wire [15:0] FP16MAC_io_c; // @[Unit.scala 422:23]
  wire [15:0] FP16MAC_io_out; // @[Unit.scala 422:23]
  reg [15:0] register_0; // @[Unit.scala 419:25]
  reg [15:0] register_1; // @[Unit.scala 419:25]
  reg [15:0] register_2; // @[Unit.scala 419:25]
  reg [15:0] register_3; // @[Unit.scala 419:25]
  reg [15:0] register_4; // @[Unit.scala 419:25]
  reg [15:0] register_5; // @[Unit.scala 419:25]
  reg [15:0] register_6; // @[Unit.scala 419:25]
  reg [15:0] register_7; // @[Unit.scala 419:25]
  reg [15:0] register_8; // @[Unit.scala 419:25]
  reg [15:0] register_9; // @[Unit.scala 419:25]
  reg [15:0] register_10; // @[Unit.scala 419:25]
  reg [15:0] register_11; // @[Unit.scala 419:25]
  reg [15:0] register_12; // @[Unit.scala 419:25]
  reg [15:0] register_13; // @[Unit.scala 419:25]
  reg [15:0] register_14; // @[Unit.scala 419:25]
  reg [15:0] register_15; // @[Unit.scala 419:25]
  reg [15:0] register_16; // @[Unit.scala 419:25]
  reg [15:0] register_17; // @[Unit.scala 419:25]
  reg [15:0] register_18; // @[Unit.scala 419:25]
  reg [15:0] register_19; // @[Unit.scala 419:25]
  reg [15:0] register_20; // @[Unit.scala 419:25]
  reg [15:0] register_21; // @[Unit.scala 419:25]
  reg [15:0] register_22; // @[Unit.scala 419:25]
  reg [15:0] register_23; // @[Unit.scala 419:25]
  reg [15:0] register_24; // @[Unit.scala 419:25]
  reg [15:0] register_25; // @[Unit.scala 419:25]
  reg [15:0] register_26; // @[Unit.scala 419:25]
  reg [15:0] register_27; // @[Unit.scala 419:25]
  reg [15:0] register_28; // @[Unit.scala 419:25]
  reg [15:0] register_29; // @[Unit.scala 419:25]
  reg [15:0] register_30; // @[Unit.scala 419:25]
  reg [15:0] register_31; // @[Unit.scala 419:25]
  reg [15:0] register_32; // @[Unit.scala 419:25]
  reg [15:0] register_33; // @[Unit.scala 419:25]
  reg [15:0] register_34; // @[Unit.scala 419:25]
  reg [15:0] register_35; // @[Unit.scala 419:25]
  reg [15:0] register_36; // @[Unit.scala 419:25]
  reg [15:0] register_37; // @[Unit.scala 419:25]
  reg [15:0] register_38; // @[Unit.scala 419:25]
  reg [15:0] register_39; // @[Unit.scala 419:25]
  reg [15:0] register_40; // @[Unit.scala 419:25]
  reg [15:0] register_41; // @[Unit.scala 419:25]
  reg [15:0] register_42; // @[Unit.scala 419:25]
  reg [15:0] register_43; // @[Unit.scala 419:25]
  reg [15:0] register_44; // @[Unit.scala 419:25]
  reg [15:0] register_45; // @[Unit.scala 419:25]
  reg [15:0] register_46; // @[Unit.scala 419:25]
  reg [15:0] register_47; // @[Unit.scala 419:25]
  reg [15:0] register_48; // @[Unit.scala 419:25]
  reg [15:0] register_49; // @[Unit.scala 419:25]
  reg [15:0] register_50; // @[Unit.scala 419:25]
  reg [15:0] register_51; // @[Unit.scala 419:25]
  reg [15:0] register_52; // @[Unit.scala 419:25]
  reg [15:0] register_53; // @[Unit.scala 419:25]
  reg [15:0] register_54; // @[Unit.scala 419:25]
  reg [15:0] register_55; // @[Unit.scala 419:25]
  reg [15:0] register_56; // @[Unit.scala 419:25]
  reg [15:0] register_57; // @[Unit.scala 419:25]
  reg [15:0] register_58; // @[Unit.scala 419:25]
  reg [15:0] register_59; // @[Unit.scala 419:25]
  reg [15:0] register_60; // @[Unit.scala 419:25]
  reg [15:0] register_61; // @[Unit.scala 419:25]
  reg [15:0] register_62; // @[Unit.scala 419:25]
  reg [15:0] register_63; // @[Unit.scala 419:25]
  wire [15:0] _GEN_3328 = io_to_PE_control == 3'h5 ? register_60 : 16'h0; // @[Unit.scala 453:38 Unit.scala 455:19 Unit.scala 463:21]
  wire [15:0] _GEN_3329 = io_to_PE_control == 3'h5 ? register_61 : 16'h0; // @[Unit.scala 453:38 Unit.scala 455:19 Unit.scala 463:21]
  wire [15:0] _GEN_3330 = io_to_PE_control == 3'h5 ? register_62 : 16'h0; // @[Unit.scala 453:38 Unit.scala 455:19 Unit.scala 463:21]
  wire [15:0] _GEN_3331 = io_to_PE_control == 3'h5 ? register_63 : 16'h0; // @[Unit.scala 453:38 Unit.scala 455:19 Unit.scala 463:21]
  wire [15:0] _GEN_3333 = io_to_PE_control == 3'h4 ? register_48 : _GEN_3328; // @[Unit.scala 448:38 Unit.scala 450:19]
  wire [15:0] _GEN_3334 = io_to_PE_control == 3'h4 ? register_49 : _GEN_3329; // @[Unit.scala 448:38 Unit.scala 450:19]
  wire [15:0] _GEN_3335 = io_to_PE_control == 3'h4 ? register_50 : _GEN_3330; // @[Unit.scala 448:38 Unit.scala 450:19]
  wire [15:0] _GEN_3336 = io_to_PE_control == 3'h4 ? register_51 : _GEN_3331; // @[Unit.scala 448:38 Unit.scala 450:19]
  wire [15:0] _GEN_3337 = io_to_PE_control == 3'h4 ? register_52 : 16'h0; // @[Unit.scala 448:38 Unit.scala 450:19]
  wire [15:0] _GEN_3338 = io_to_PE_control == 3'h4 ? register_53 : 16'h0; // @[Unit.scala 448:38 Unit.scala 450:19]
  wire [15:0] _GEN_3339 = io_to_PE_control == 3'h4 ? register_54 : 16'h0; // @[Unit.scala 448:38 Unit.scala 450:19]
  wire [15:0] _GEN_3340 = io_to_PE_control == 3'h4 ? register_55 : 16'h0; // @[Unit.scala 448:38 Unit.scala 450:19]
  wire [15:0] _GEN_3341 = io_to_PE_control == 3'h4 ? register_56 : 16'h0; // @[Unit.scala 448:38 Unit.scala 450:19]
  wire [15:0] _GEN_3342 = io_to_PE_control == 3'h4 ? register_57 : 16'h0; // @[Unit.scala 448:38 Unit.scala 450:19]
  wire [15:0] _GEN_3343 = io_to_PE_control == 3'h4 ? register_58 : 16'h0; // @[Unit.scala 448:38 Unit.scala 450:19]
  wire [15:0] _GEN_3344 = io_to_PE_control == 3'h4 ? register_59 : 16'h0; // @[Unit.scala 448:38 Unit.scala 450:19]
  wire [15:0] _GEN_3345 = io_to_PE_control == 3'h3 ? register_36 : _GEN_3333; // @[Unit.scala 443:38 Unit.scala 445:19]
  wire [15:0] _GEN_3346 = io_to_PE_control == 3'h3 ? register_37 : _GEN_3334; // @[Unit.scala 443:38 Unit.scala 445:19]
  wire [15:0] _GEN_3347 = io_to_PE_control == 3'h3 ? register_38 : _GEN_3335; // @[Unit.scala 443:38 Unit.scala 445:19]
  wire [15:0] _GEN_3348 = io_to_PE_control == 3'h3 ? register_39 : _GEN_3336; // @[Unit.scala 443:38 Unit.scala 445:19]
  wire [15:0] _GEN_3349 = io_to_PE_control == 3'h3 ? register_40 : _GEN_3337; // @[Unit.scala 443:38 Unit.scala 445:19]
  wire [15:0] _GEN_3350 = io_to_PE_control == 3'h3 ? register_41 : _GEN_3338; // @[Unit.scala 443:38 Unit.scala 445:19]
  wire [15:0] _GEN_3351 = io_to_PE_control == 3'h3 ? register_42 : _GEN_3339; // @[Unit.scala 443:38 Unit.scala 445:19]
  wire [15:0] _GEN_3352 = io_to_PE_control == 3'h3 ? register_43 : _GEN_3340; // @[Unit.scala 443:38 Unit.scala 445:19]
  wire [15:0] _GEN_3353 = io_to_PE_control == 3'h3 ? register_44 : _GEN_3341; // @[Unit.scala 443:38 Unit.scala 445:19]
  wire [15:0] _GEN_3354 = io_to_PE_control == 3'h3 ? register_45 : _GEN_3342; // @[Unit.scala 443:38 Unit.scala 445:19]
  wire [15:0] _GEN_3355 = io_to_PE_control == 3'h3 ? register_46 : _GEN_3343; // @[Unit.scala 443:38 Unit.scala 445:19]
  wire [15:0] _GEN_3356 = io_to_PE_control == 3'h3 ? register_47 : _GEN_3344; // @[Unit.scala 443:38 Unit.scala 445:19]
  wire [15:0] _GEN_3357 = io_to_PE_control == 3'h2 ? register_24 : _GEN_3345; // @[Unit.scala 438:38 Unit.scala 440:19]
  wire [15:0] _GEN_3358 = io_to_PE_control == 3'h2 ? register_25 : _GEN_3346; // @[Unit.scala 438:38 Unit.scala 440:19]
  wire [15:0] _GEN_3359 = io_to_PE_control == 3'h2 ? register_26 : _GEN_3347; // @[Unit.scala 438:38 Unit.scala 440:19]
  wire [15:0] _GEN_3360 = io_to_PE_control == 3'h2 ? register_27 : _GEN_3348; // @[Unit.scala 438:38 Unit.scala 440:19]
  wire [15:0] _GEN_3361 = io_to_PE_control == 3'h2 ? register_28 : _GEN_3349; // @[Unit.scala 438:38 Unit.scala 440:19]
  wire [15:0] _GEN_3362 = io_to_PE_control == 3'h2 ? register_29 : _GEN_3350; // @[Unit.scala 438:38 Unit.scala 440:19]
  wire [15:0] _GEN_3363 = io_to_PE_control == 3'h2 ? register_30 : _GEN_3351; // @[Unit.scala 438:38 Unit.scala 440:19]
  wire [15:0] _GEN_3364 = io_to_PE_control == 3'h2 ? register_31 : _GEN_3352; // @[Unit.scala 438:38 Unit.scala 440:19]
  wire [15:0] _GEN_3365 = io_to_PE_control == 3'h2 ? register_0 : _GEN_3353; // @[Unit.scala 438:38 Unit.scala 440:19]
  wire [15:0] _GEN_3366 = io_to_PE_control == 3'h2 ? register_1 : _GEN_3354; // @[Unit.scala 438:38 Unit.scala 440:19]
  wire [15:0] _GEN_3367 = io_to_PE_control == 3'h2 ? register_2 : _GEN_3355; // @[Unit.scala 438:38 Unit.scala 440:19]
  wire [15:0] _GEN_3368 = io_to_PE_control == 3'h2 ? register_3 : _GEN_3356; // @[Unit.scala 438:38 Unit.scala 440:19]
  wire [15:0] _GEN_3369 = io_to_PE_control == 3'h1 ? register_12 : _GEN_3357; // @[Unit.scala 433:38 Unit.scala 435:19]
  wire [15:0] _GEN_3370 = io_to_PE_control == 3'h1 ? register_13 : _GEN_3358; // @[Unit.scala 433:38 Unit.scala 435:19]
  wire [15:0] _GEN_3371 = io_to_PE_control == 3'h1 ? register_14 : _GEN_3359; // @[Unit.scala 433:38 Unit.scala 435:19]
  wire [15:0] _GEN_3372 = io_to_PE_control == 3'h1 ? register_15 : _GEN_3360; // @[Unit.scala 433:38 Unit.scala 435:19]
  wire [15:0] _GEN_3373 = io_to_PE_control == 3'h1 ? register_0 : _GEN_3361; // @[Unit.scala 433:38 Unit.scala 435:19]
  wire [15:0] _GEN_3374 = io_to_PE_control == 3'h1 ? register_1 : _GEN_3362; // @[Unit.scala 433:38 Unit.scala 435:19]
  wire [15:0] _GEN_3375 = io_to_PE_control == 3'h1 ? register_2 : _GEN_3363; // @[Unit.scala 433:38 Unit.scala 435:19]
  wire [15:0] _GEN_3376 = io_to_PE_control == 3'h1 ? register_3 : _GEN_3364; // @[Unit.scala 433:38 Unit.scala 435:19]
  wire [15:0] _GEN_3377 = io_to_PE_control == 3'h1 ? register_4 : _GEN_3365; // @[Unit.scala 433:38 Unit.scala 435:19]
  wire [15:0] _GEN_3378 = io_to_PE_control == 3'h1 ? register_5 : _GEN_3366; // @[Unit.scala 433:38 Unit.scala 435:19]
  wire [15:0] _GEN_3379 = io_to_PE_control == 3'h1 ? register_6 : _GEN_3367; // @[Unit.scala 433:38 Unit.scala 435:19]
  wire [15:0] _GEN_3380 = io_to_PE_control == 3'h1 ? register_7 : _GEN_3368; // @[Unit.scala 433:38 Unit.scala 435:19]
  wire [15:0] _GEN_3458 = 6'h1 == io_wrAddr ? register_1 : register_0; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3459 = 6'h2 == io_wrAddr ? register_2 : _GEN_3458; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3460 = 6'h3 == io_wrAddr ? register_3 : _GEN_3459; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3461 = 6'h4 == io_wrAddr ? register_4 : _GEN_3460; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3462 = 6'h5 == io_wrAddr ? register_5 : _GEN_3461; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3463 = 6'h6 == io_wrAddr ? register_6 : _GEN_3462; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3464 = 6'h7 == io_wrAddr ? register_7 : _GEN_3463; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3465 = 6'h8 == io_wrAddr ? register_8 : _GEN_3464; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3466 = 6'h9 == io_wrAddr ? register_9 : _GEN_3465; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3467 = 6'ha == io_wrAddr ? register_10 : _GEN_3466; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3468 = 6'hb == io_wrAddr ? register_11 : _GEN_3467; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3469 = 6'hc == io_wrAddr ? register_12 : _GEN_3468; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3470 = 6'hd == io_wrAddr ? register_13 : _GEN_3469; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3471 = 6'he == io_wrAddr ? register_14 : _GEN_3470; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3472 = 6'hf == io_wrAddr ? register_15 : _GEN_3471; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3473 = 6'h10 == io_wrAddr ? register_16 : _GEN_3472; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3474 = 6'h11 == io_wrAddr ? register_17 : _GEN_3473; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3475 = 6'h12 == io_wrAddr ? register_18 : _GEN_3474; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3476 = 6'h13 == io_wrAddr ? register_19 : _GEN_3475; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3477 = 6'h14 == io_wrAddr ? register_20 : _GEN_3476; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3478 = 6'h15 == io_wrAddr ? register_21 : _GEN_3477; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3479 = 6'h16 == io_wrAddr ? register_22 : _GEN_3478; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3480 = 6'h17 == io_wrAddr ? register_23 : _GEN_3479; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3481 = 6'h18 == io_wrAddr ? register_24 : _GEN_3480; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3482 = 6'h19 == io_wrAddr ? register_25 : _GEN_3481; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3483 = 6'h1a == io_wrAddr ? register_26 : _GEN_3482; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3484 = 6'h1b == io_wrAddr ? register_27 : _GEN_3483; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3485 = 6'h1c == io_wrAddr ? register_28 : _GEN_3484; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3486 = 6'h1d == io_wrAddr ? register_29 : _GEN_3485; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3487 = 6'h1e == io_wrAddr ? register_30 : _GEN_3486; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3488 = 6'h1f == io_wrAddr ? register_31 : _GEN_3487; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3489 = 6'h20 == io_wrAddr ? register_32 : _GEN_3488; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3490 = 6'h21 == io_wrAddr ? register_33 : _GEN_3489; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3491 = 6'h22 == io_wrAddr ? register_34 : _GEN_3490; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3492 = 6'h23 == io_wrAddr ? register_35 : _GEN_3491; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3493 = 6'h24 == io_wrAddr ? register_36 : _GEN_3492; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3494 = 6'h25 == io_wrAddr ? register_37 : _GEN_3493; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3495 = 6'h26 == io_wrAddr ? register_38 : _GEN_3494; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3496 = 6'h27 == io_wrAddr ? register_39 : _GEN_3495; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3497 = 6'h28 == io_wrAddr ? register_40 : _GEN_3496; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3498 = 6'h29 == io_wrAddr ? register_41 : _GEN_3497; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3499 = 6'h2a == io_wrAddr ? register_42 : _GEN_3498; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3500 = 6'h2b == io_wrAddr ? register_43 : _GEN_3499; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3501 = 6'h2c == io_wrAddr ? register_44 : _GEN_3500; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3502 = 6'h2d == io_wrAddr ? register_45 : _GEN_3501; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3503 = 6'h2e == io_wrAddr ? register_46 : _GEN_3502; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3504 = 6'h2f == io_wrAddr ? register_47 : _GEN_3503; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3505 = 6'h30 == io_wrAddr ? register_48 : _GEN_3504; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3506 = 6'h31 == io_wrAddr ? register_49 : _GEN_3505; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3507 = 6'h32 == io_wrAddr ? register_50 : _GEN_3506; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3508 = 6'h33 == io_wrAddr ? register_51 : _GEN_3507; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3509 = 6'h34 == io_wrAddr ? register_52 : _GEN_3508; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3510 = 6'h35 == io_wrAddr ? register_53 : _GEN_3509; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3511 = 6'h36 == io_wrAddr ? register_54 : _GEN_3510; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3512 = 6'h37 == io_wrAddr ? register_55 : _GEN_3511; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3513 = 6'h38 == io_wrAddr ? register_56 : _GEN_3512; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3514 = 6'h39 == io_wrAddr ? register_57 : _GEN_3513; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3515 = 6'h3a == io_wrAddr ? register_58 : _GEN_3514; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3516 = 6'h3b == io_wrAddr ? register_59 : _GEN_3515; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3517 = 6'h3c == io_wrAddr ? register_60 : _GEN_3516; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3518 = 6'h3d == io_wrAddr ? register_61 : _GEN_3517; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3519 = 6'h3e == io_wrAddr ? register_62 : _GEN_3518; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _GEN_3520 = 6'h3f == io_wrAddr ? register_63 : _GEN_3519; // @[Unit.scala 473:18 Unit.scala 473:18]
  wire [15:0] _register_io_wrAddr_0 = FP16MAC_io_out; // @[Unit.scala 474:25 Unit.scala 474:25]
  wire [13:0] _GEN_3586 = io_wrEna ? 14'h3c00 : 14'h0; // @[Unit.scala 470:18 Unit.scala 472:18 Unit.scala 478:20]
  FP16MulAdder FP16MAC ( // @[Unit.scala 422:23]
    .io_a(FP16MAC_io_a),
    .io_b(FP16MAC_io_b),
    .io_c(FP16MAC_io_c),
    .io_out(FP16MAC_io_out)
  );
  assign io_to_PE_0 = io_to_PE_control == 3'h0 ? register_0 : _GEN_3369; // @[Unit.scala 428:33 Unit.scala 430:19]
  assign io_to_PE_1 = io_to_PE_control == 3'h0 ? register_1 : _GEN_3370; // @[Unit.scala 428:33 Unit.scala 430:19]
  assign io_to_PE_2 = io_to_PE_control == 3'h0 ? register_2 : _GEN_3371; // @[Unit.scala 428:33 Unit.scala 430:19]
  assign io_to_PE_3 = io_to_PE_control == 3'h0 ? register_3 : _GEN_3372; // @[Unit.scala 428:33 Unit.scala 430:19]
  assign io_to_PE_4 = io_to_PE_control == 3'h0 ? register_4 : _GEN_3373; // @[Unit.scala 428:33 Unit.scala 430:19]
  assign io_to_PE_5 = io_to_PE_control == 3'h0 ? register_5 : _GEN_3374; // @[Unit.scala 428:33 Unit.scala 430:19]
  assign io_to_PE_6 = io_to_PE_control == 3'h0 ? register_6 : _GEN_3375; // @[Unit.scala 428:33 Unit.scala 430:19]
  assign io_to_PE_7 = io_to_PE_control == 3'h0 ? register_7 : _GEN_3376; // @[Unit.scala 428:33 Unit.scala 430:19]
  assign io_to_PE_8 = io_to_PE_control == 3'h0 ? register_8 : _GEN_3377; // @[Unit.scala 428:33 Unit.scala 430:19]
  assign io_to_PE_9 = io_to_PE_control == 3'h0 ? register_9 : _GEN_3378; // @[Unit.scala 428:33 Unit.scala 430:19]
  assign io_to_PE_10 = io_to_PE_control == 3'h0 ? register_10 : _GEN_3379; // @[Unit.scala 428:33 Unit.scala 430:19]
  assign io_to_PE_11 = io_to_PE_control == 3'h0 ? register_11 : _GEN_3380; // @[Unit.scala 428:33 Unit.scala 430:19]
  assign io_rdData = register_0; // @[Unit.scala 468:13 Unit.scala 468:13]
  assign FP16MAC_io_a = io_wrEna ? io_wrData : 16'h0; // @[Unit.scala 470:18 Unit.scala 471:18 Unit.scala 477:20]
  assign FP16MAC_io_b = {{2'd0}, _GEN_3586}; // @[Unit.scala 470:18 Unit.scala 472:18 Unit.scala 478:20]
  assign FP16MAC_io_c = io_wrEna ? _GEN_3520 : 16'h0; // @[Unit.scala 470:18 Unit.scala 473:18 Unit.scala 479:20]
  always @(posedge clock) begin
    if (reset) begin // @[Unit.scala 419:25]
      register_0 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h0 == io_wrAddr) begin // @[Unit.scala 474:25]
        register_0 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_1 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h1 == io_wrAddr) begin // @[Unit.scala 474:25]
        register_1 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_2 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h2 == io_wrAddr) begin // @[Unit.scala 474:25]
        register_2 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_3 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h3 == io_wrAddr) begin // @[Unit.scala 474:25]
        register_3 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_4 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h4 == io_wrAddr) begin // @[Unit.scala 474:25]
        register_4 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_5 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h5 == io_wrAddr) begin // @[Unit.scala 474:25]
        register_5 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_6 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h6 == io_wrAddr) begin // @[Unit.scala 474:25]
        register_6 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_7 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h7 == io_wrAddr) begin // @[Unit.scala 474:25]
        register_7 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_8 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h8 == io_wrAddr) begin // @[Unit.scala 474:25]
        register_8 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_9 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h9 == io_wrAddr) begin // @[Unit.scala 474:25]
        register_9 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_10 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'ha == io_wrAddr) begin // @[Unit.scala 474:25]
        register_10 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_11 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'hb == io_wrAddr) begin // @[Unit.scala 474:25]
        register_11 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_12 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'hc == io_wrAddr) begin // @[Unit.scala 474:25]
        register_12 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_13 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'hd == io_wrAddr) begin // @[Unit.scala 474:25]
        register_13 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_14 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'he == io_wrAddr) begin // @[Unit.scala 474:25]
        register_14 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_15 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'hf == io_wrAddr) begin // @[Unit.scala 474:25]
        register_15 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_16 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h10 == io_wrAddr) begin // @[Unit.scala 474:25]
        register_16 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_17 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h11 == io_wrAddr) begin // @[Unit.scala 474:25]
        register_17 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_18 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h12 == io_wrAddr) begin // @[Unit.scala 474:25]
        register_18 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_19 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h13 == io_wrAddr) begin // @[Unit.scala 474:25]
        register_19 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_20 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h14 == io_wrAddr) begin // @[Unit.scala 474:25]
        register_20 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_21 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h15 == io_wrAddr) begin // @[Unit.scala 474:25]
        register_21 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_22 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h16 == io_wrAddr) begin // @[Unit.scala 474:25]
        register_22 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_23 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h17 == io_wrAddr) begin // @[Unit.scala 474:25]
        register_23 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_24 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h18 == io_wrAddr) begin // @[Unit.scala 474:25]
        register_24 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_25 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h19 == io_wrAddr) begin // @[Unit.scala 474:25]
        register_25 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_26 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h1a == io_wrAddr) begin // @[Unit.scala 474:25]
        register_26 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_27 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h1b == io_wrAddr) begin // @[Unit.scala 474:25]
        register_27 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_28 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h1c == io_wrAddr) begin // @[Unit.scala 474:25]
        register_28 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_29 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h1d == io_wrAddr) begin // @[Unit.scala 474:25]
        register_29 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_30 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h1e == io_wrAddr) begin // @[Unit.scala 474:25]
        register_30 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_31 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h1f == io_wrAddr) begin // @[Unit.scala 474:25]
        register_31 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_32 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h20 == io_wrAddr) begin // @[Unit.scala 474:25]
        register_32 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_33 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h21 == io_wrAddr) begin // @[Unit.scala 474:25]
        register_33 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_34 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h22 == io_wrAddr) begin // @[Unit.scala 474:25]
        register_34 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_35 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h23 == io_wrAddr) begin // @[Unit.scala 474:25]
        register_35 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_36 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h24 == io_wrAddr) begin // @[Unit.scala 474:25]
        register_36 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_37 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h25 == io_wrAddr) begin // @[Unit.scala 474:25]
        register_37 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_38 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h26 == io_wrAddr) begin // @[Unit.scala 474:25]
        register_38 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_39 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h27 == io_wrAddr) begin // @[Unit.scala 474:25]
        register_39 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_40 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h28 == io_wrAddr) begin // @[Unit.scala 474:25]
        register_40 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_41 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h29 == io_wrAddr) begin // @[Unit.scala 474:25]
        register_41 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_42 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h2a == io_wrAddr) begin // @[Unit.scala 474:25]
        register_42 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_43 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h2b == io_wrAddr) begin // @[Unit.scala 474:25]
        register_43 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_44 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h2c == io_wrAddr) begin // @[Unit.scala 474:25]
        register_44 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_45 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h2d == io_wrAddr) begin // @[Unit.scala 474:25]
        register_45 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_46 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h2e == io_wrAddr) begin // @[Unit.scala 474:25]
        register_46 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_47 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h2f == io_wrAddr) begin // @[Unit.scala 474:25]
        register_47 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_48 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h30 == io_wrAddr) begin // @[Unit.scala 474:25]
        register_48 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_49 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h31 == io_wrAddr) begin // @[Unit.scala 474:25]
        register_49 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_50 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h32 == io_wrAddr) begin // @[Unit.scala 474:25]
        register_50 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_51 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h33 == io_wrAddr) begin // @[Unit.scala 474:25]
        register_51 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_52 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h34 == io_wrAddr) begin // @[Unit.scala 474:25]
        register_52 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_53 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h35 == io_wrAddr) begin // @[Unit.scala 474:25]
        register_53 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_54 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h36 == io_wrAddr) begin // @[Unit.scala 474:25]
        register_54 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_55 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h37 == io_wrAddr) begin // @[Unit.scala 474:25]
        register_55 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_56 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h38 == io_wrAddr) begin // @[Unit.scala 474:25]
        register_56 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_57 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h39 == io_wrAddr) begin // @[Unit.scala 474:25]
        register_57 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_58 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h3a == io_wrAddr) begin // @[Unit.scala 474:25]
        register_58 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_59 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h3b == io_wrAddr) begin // @[Unit.scala 474:25]
        register_59 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_60 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h3c == io_wrAddr) begin // @[Unit.scala 474:25]
        register_60 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_61 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h3d == io_wrAddr) begin // @[Unit.scala 474:25]
        register_61 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_62 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h3e == io_wrAddr) begin // @[Unit.scala 474:25]
        register_62 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
    if (reset) begin // @[Unit.scala 419:25]
      register_63 <= 16'h0; // @[Unit.scala 419:25]
    end else if (io_wrEna) begin // @[Unit.scala 470:18]
      if (6'h3f == io_wrAddr) begin // @[Unit.scala 474:25]
        register_63 <= _register_io_wrAddr_0; // @[Unit.scala 474:25]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  register_0 = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  register_1 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  register_2 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  register_3 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  register_4 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  register_5 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  register_6 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  register_7 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  register_8 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  register_9 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  register_10 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  register_11 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  register_12 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  register_13 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  register_14 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  register_15 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  register_16 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  register_17 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  register_18 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  register_19 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  register_20 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  register_21 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  register_22 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  register_23 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  register_24 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  register_25 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  register_26 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  register_27 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  register_28 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  register_29 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  register_30 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  register_31 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  register_32 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  register_33 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  register_34 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  register_35 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  register_36 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  register_37 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  register_38 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  register_39 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  register_40 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  register_41 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  register_42 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  register_43 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  register_44 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  register_45 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  register_46 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  register_47 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  register_48 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  register_49 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  register_50 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  register_51 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  register_52 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  register_53 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  register_54 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  register_55 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  register_56 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  register_57 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  register_58 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  register_59 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  register_60 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  register_61 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  register_62 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  register_63 = _RAND_63[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module tanh_Unit(
  input  [15:0] io_input,
  output [15:0] io_output
);
  wire [15:0] FP16MAC_io_a; // @[Unit.scala 286:23]
  wire [15:0] FP16MAC_io_b; // @[Unit.scala 286:23]
  wire [15:0] FP16MAC_io_c; // @[Unit.scala 286:23]
  wire [15:0] FP16MAC_io_out; // @[Unit.scala 286:23]
  wire  _T_39 = ~io_input[15]; // @[Unit.scala 333:36]
  wire [15:0] _GEN_0 = _T_39 & io_input > 16'h4500 & io_input <= 16'h4600 ? io_input : 16'h0; // @[Unit.scala 363:98 Unit.scala 364:20 Unit.scala 371:20]
  wire [12:0] _GEN_1 = _T_39 & io_input > 16'h4500 & io_input <= 16'h4600 ? 13'h1c4d : 13'h0; // @[Unit.scala 363:98 Unit.scala 365:20 Unit.scala 372:20]
  wire [13:0] _GEN_2 = _T_39 & io_input > 16'h4500 & io_input <= 16'h4600 ? 14'h3bc8 : 14'h0; // @[Unit.scala 363:98 Unit.scala 366:20 Unit.scala 373:20]
  wire [15:0] _GEN_3 = _T_39 & io_input > 16'h4500 & io_input <= 16'h4600 ? FP16MAC_io_out : 16'h3c00; // @[Unit.scala 363:98 Unit.scala 367:17 Unit.scala 370:17]
  wire [15:0] _GEN_4 = _T_39 & io_input > 16'h4400 & io_input <= 16'h4500 ? io_input : _GEN_0; // @[Unit.scala 357:98 Unit.scala 358:20]
  wire [13:0] _GEN_5 = _T_39 & io_input > 16'h4400 & io_input <= 16'h4500 ? 14'h21ae : {{1'd0}, _GEN_1}; // @[Unit.scala 357:98 Unit.scala 359:20]
  wire [13:0] _GEN_6 = _T_39 & io_input > 16'h4400 & io_input <= 16'h4500 ? 14'h3b82 : _GEN_2; // @[Unit.scala 357:98 Unit.scala 360:20]
  wire [15:0] _GEN_7 = _T_39 & io_input > 16'h4400 & io_input <= 16'h4500 ? FP16MAC_io_out : _GEN_3; // @[Unit.scala 357:98 Unit.scala 361:17]
  wire [15:0] _GEN_8 = _T_39 & io_input > 16'h4200 & io_input <= 16'h4400 ? io_input : _GEN_4; // @[Unit.scala 351:98 Unit.scala 352:20]
  wire [13:0] _GEN_9 = _T_39 & io_input > 16'h4200 & io_input <= 16'h4400 ? 14'h2773 : _GEN_5; // @[Unit.scala 351:98 Unit.scala 353:20]
  wire [13:0] _GEN_10 = _T_39 & io_input > 16'h4200 & io_input <= 16'h4400 ? 14'h3af1 : _GEN_6; // @[Unit.scala 351:98 Unit.scala 354:20]
  wire [15:0] _GEN_11 = _T_39 & io_input > 16'h4200 & io_input <= 16'h4400 ? FP16MAC_io_out : _GEN_7; // @[Unit.scala 351:98 Unit.scala 355:17]
  wire [15:0] _GEN_12 = _T_39 & io_input > 16'h4000 & io_input <= 16'h4200 ? io_input : _GEN_8; // @[Unit.scala 345:98 Unit.scala 346:20]
  wire [13:0] _GEN_13 = _T_39 & io_input > 16'h4000 & io_input <= 16'h4200 ? 14'h2c8c : _GEN_9; // @[Unit.scala 345:98 Unit.scala 347:20]
  wire [13:0] _GEN_14 = _T_39 & io_input > 16'h4000 & io_input <= 16'h4200 ? 14'h39f3 : _GEN_10; // @[Unit.scala 345:98 Unit.scala 348:20]
  wire [15:0] _GEN_15 = _T_39 & io_input > 16'h4000 & io_input <= 16'h4200 ? FP16MAC_io_out : _GEN_11; // @[Unit.scala 345:98 Unit.scala 349:17]
  wire [15:0] _GEN_16 = _T_39 & io_input > 16'h3c00 & io_input <= 16'h4000 ? io_input : _GEN_12; // @[Unit.scala 339:98 Unit.scala 340:20]
  wire [13:0] _GEN_17 = _T_39 & io_input > 16'h3c00 & io_input <= 16'h4000 ? 14'h30c8 : _GEN_13; // @[Unit.scala 339:98 Unit.scala 341:20]
  wire [13:0] _GEN_18 = _T_39 & io_input > 16'h3c00 & io_input <= 16'h4000 ? 14'h38b6 : _GEN_14; // @[Unit.scala 339:98 Unit.scala 342:20]
  wire [15:0] _GEN_19 = _T_39 & io_input > 16'h3c00 & io_input <= 16'h4000 ? FP16MAC_io_out : _GEN_15; // @[Unit.scala 339:98 Unit.scala 343:17]
  wire [15:0] _GEN_20 = ~io_input[15] & io_input <= 16'h3c00 ? io_input : _GEN_16; // @[Unit.scala 333:93 Unit.scala 334:20]
  wire [13:0] _GEN_21 = ~io_input[15] & io_input <= 16'h3c00 ? 14'h3371 : _GEN_17; // @[Unit.scala 333:93 Unit.scala 335:20]
  wire [13:0] _GEN_22 = ~io_input[15] & io_input <= 16'h3c00 ? 14'h3807 : _GEN_18; // @[Unit.scala 333:93 Unit.scala 336:20]
  wire [15:0] _GEN_23 = ~io_input[15] & io_input <= 16'h3c00 ? FP16MAC_io_out : _GEN_19; // @[Unit.scala 333:93 Unit.scala 337:17]
  wire [15:0] _GEN_24 = io_input[15] & io_input < 16'hbc00 ? io_input : _GEN_20; // @[Unit.scala 327:71 Unit.scala 328:20]
  wire [13:0] _GEN_25 = io_input[15] & io_input < 16'hbc00 ? 14'h3371 : _GEN_21; // @[Unit.scala 327:71 Unit.scala 329:20]
  wire [13:0] _GEN_26 = io_input[15] & io_input < 16'hbc00 ? 14'h37f0 : _GEN_22; // @[Unit.scala 327:71 Unit.scala 330:20]
  wire [15:0] _GEN_27 = io_input[15] & io_input < 16'hbc00 ? FP16MAC_io_out : _GEN_23; // @[Unit.scala 327:71 Unit.scala 331:17]
  wire [15:0] _GEN_28 = io_input[15] & io_input < 16'hc000 & io_input >= 16'hbc00 ? io_input : _GEN_24; // @[Unit.scala 321:98 Unit.scala 322:20]
  wire [13:0] _GEN_29 = io_input[15] & io_input < 16'hc000 & io_input >= 16'hbc00 ? 14'h30c8 : _GEN_25; // @[Unit.scala 321:98 Unit.scala 323:20]
  wire [13:0] _GEN_30 = io_input[15] & io_input < 16'hc000 & io_input >= 16'hbc00 ? 14'h3692 : _GEN_26; // @[Unit.scala 321:98 Unit.scala 324:20]
  wire [15:0] _GEN_31 = io_input[15] & io_input < 16'hc000 & io_input >= 16'hbc00 ? FP16MAC_io_out : _GEN_27; // @[Unit.scala 321:98 Unit.scala 325:17]
  wire [15:0] _GEN_32 = io_input[15] & io_input < 16'hc200 & io_input >= 16'hc000 ? io_input : _GEN_28; // @[Unit.scala 315:98 Unit.scala 316:20]
  wire [13:0] _GEN_33 = io_input[15] & io_input < 16'hc200 & io_input >= 16'hc000 ? 14'h2c8c : _GEN_29; // @[Unit.scala 315:98 Unit.scala 317:20]
  wire [13:0] _GEN_34 = io_input[15] & io_input < 16'hc200 & io_input >= 16'hc000 ? 14'h3419 : _GEN_30; // @[Unit.scala 315:98 Unit.scala 318:20]
  wire [15:0] _GEN_35 = io_input[15] & io_input < 16'hc200 & io_input >= 16'hc000 ? FP16MAC_io_out : _GEN_31; // @[Unit.scala 315:98 Unit.scala 319:17]
  wire [15:0] _GEN_36 = io_input[15] & io_input < 16'hc400 & io_input >= 16'hc200 ? io_input : _GEN_32; // @[Unit.scala 309:98 Unit.scala 310:20]
  wire [13:0] _GEN_37 = io_input[15] & io_input < 16'hc400 & io_input >= 16'hc200 ? 14'h2773 : _GEN_33; // @[Unit.scala 309:98 Unit.scala 311:20]
  wire [13:0] _GEN_38 = io_input[15] & io_input < 16'hc400 & io_input >= 16'hc200 ? 14'h303a : _GEN_34; // @[Unit.scala 309:98 Unit.scala 312:20]
  wire [15:0] _GEN_39 = io_input[15] & io_input < 16'hc400 & io_input >= 16'hc200 ? FP16MAC_io_out : _GEN_35; // @[Unit.scala 309:98 Unit.scala 313:17]
  wire [15:0] _GEN_40 = io_input[15] & io_input < 16'hc500 & io_input >= 16'hc400 ? io_input : _GEN_36; // @[Unit.scala 303:98 Unit.scala 304:20]
  wire [13:0] _GEN_41 = io_input[15] & io_input < 16'hc500 & io_input >= 16'hc400 ? 14'h21ae : _GEN_37; // @[Unit.scala 303:98 Unit.scala 305:20]
  wire [13:0] _GEN_42 = io_input[15] & io_input < 16'hc500 & io_input >= 16'hc400 ? 14'h2bdf : _GEN_38; // @[Unit.scala 303:98 Unit.scala 306:20]
  wire [15:0] _GEN_43 = io_input[15] & io_input < 16'hc500 & io_input >= 16'hc400 ? FP16MAC_io_out : _GEN_39; // @[Unit.scala 303:98 Unit.scala 307:17]
  wire [15:0] _GEN_44 = io_input[15] & io_input < 16'hc600 & io_input >= 16'hc500 ? io_input : _GEN_40; // @[Unit.scala 297:98 Unit.scala 298:20]
  wire [13:0] _GEN_45 = io_input[15] & io_input < 16'hc600 & io_input >= 16'hc500 ? 14'h1c4d : _GEN_41; // @[Unit.scala 297:98 Unit.scala 299:20]
  wire [13:0] _GEN_46 = io_input[15] & io_input < 16'hc600 & io_input >= 16'hc500 ? 14'h26f0 : _GEN_42; // @[Unit.scala 297:98 Unit.scala 300:20]
  wire [15:0] _GEN_47 = io_input[15] & io_input < 16'hc600 & io_input >= 16'hc500 ? FP16MAC_io_out : _GEN_43; // @[Unit.scala 297:98 Unit.scala 301:17]
  wire [13:0] _GEN_49 = io_input[15] & io_input >= 16'hc600 ? 14'h0 : _GEN_45; // @[Unit.scala 291:65 Unit.scala 293:18]
  wire [13:0] _GEN_50 = io_input[15] & io_input >= 16'hc600 ? 14'h0 : _GEN_46; // @[Unit.scala 291:65 Unit.scala 294:18]
  FP16MulAdder FP16MAC ( // @[Unit.scala 286:23]
    .io_a(FP16MAC_io_a),
    .io_b(FP16MAC_io_b),
    .io_c(FP16MAC_io_c),
    .io_out(FP16MAC_io_out)
  );
  assign io_output = io_input[15] & io_input >= 16'hc600 ? 16'hbc00 : _GEN_47; // @[Unit.scala 291:65 Unit.scala 295:15]
  assign FP16MAC_io_a = io_input[15] & io_input >= 16'hc600 ? 16'h0 : _GEN_44; // @[Unit.scala 291:65 Unit.scala 292:18]
  assign FP16MAC_io_b = {{2'd0}, _GEN_49}; // @[Unit.scala 291:65 Unit.scala 293:18]
  assign FP16MAC_io_c = {{2'd0}, _GEN_50}; // @[Unit.scala 291:65 Unit.scala 294:18]
endmodule
module EW_Unit(
  input         clock,
  input         reset,
  input  [15:0] io_ht_1_input,
  input  [15:0] io_Zt_input,
  input  [15:0] io_Rt_input,
  input  [15:0] io_Whxt_input,
  input  [15:0] io_Uhht_1_input,
  output [15:0] io_output
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] FP16MAC1_io_a; // @[Unit.scala 502:24]
  wire [15:0] FP16MAC1_io_b; // @[Unit.scala 502:24]
  wire [15:0] FP16MAC1_io_c; // @[Unit.scala 502:24]
  wire [15:0] FP16MAC1_io_out; // @[Unit.scala 502:24]
  wire [15:0] FP16MAC2_io_a; // @[Unit.scala 506:24]
  wire [15:0] FP16MAC2_io_b; // @[Unit.scala 506:24]
  wire [15:0] FP16MAC2_io_c; // @[Unit.scala 506:24]
  wire [15:0] FP16MAC2_io_out; // @[Unit.scala 506:24]
  wire [15:0] FP16MAC3_io_a; // @[Unit.scala 510:24]
  wire [15:0] FP16MAC3_io_b; // @[Unit.scala 510:24]
  wire [15:0] FP16MAC3_io_c; // @[Unit.scala 510:24]
  wire [15:0] FP16MAC3_io_out; // @[Unit.scala 510:24]
  wire [15:0] FP16MAC4_io_a; // @[Unit.scala 514:24]
  wire [15:0] FP16MAC4_io_b; // @[Unit.scala 514:24]
  wire [15:0] FP16MAC4_io_c; // @[Unit.scala 514:24]
  wire [15:0] FP16MAC4_io_out; // @[Unit.scala 514:24]
  wire [15:0] tanh_io_input; // @[Unit.scala 527:20]
  wire [15:0] tanh_io_output; // @[Unit.scala 527:20]
  reg [15:0] reg_before_tanh; // @[Unit.scala 493:32]
  reg [15:0] reg_Zt; // @[Unit.scala 494:30]
  reg [15:0] reg_ht_1; // @[Unit.scala 495:30]
  reg [15:0] reg_tanh; // @[Unit.scala 496:30]
  reg [15:0] reg_1_Zt; // @[Unit.scala 497:30]
  reg [15:0] reg_Zt_ht_1; // @[Unit.scala 498:30]
  reg [15:0] reg_output; // @[Unit.scala 499:30]
  wire  reg_Zt_inv_hi = ~reg_Zt[15]; // @[Unit.scala 532:24]
  wire [14:0] reg_Zt_inv_lo = reg_Zt[14:0]; // @[Unit.scala 532:49]
  FP16MulAdder FP16MAC1 ( // @[Unit.scala 502:24]
    .io_a(FP16MAC1_io_a),
    .io_b(FP16MAC1_io_b),
    .io_c(FP16MAC1_io_c),
    .io_out(FP16MAC1_io_out)
  );
  FP16MulAdder FP16MAC2 ( // @[Unit.scala 506:24]
    .io_a(FP16MAC2_io_a),
    .io_b(FP16MAC2_io_b),
    .io_c(FP16MAC2_io_c),
    .io_out(FP16MAC2_io_out)
  );
  FP16MulAdder FP16MAC3 ( // @[Unit.scala 510:24]
    .io_a(FP16MAC3_io_a),
    .io_b(FP16MAC3_io_b),
    .io_c(FP16MAC3_io_c),
    .io_out(FP16MAC3_io_out)
  );
  FP16MulAdder FP16MAC4 ( // @[Unit.scala 514:24]
    .io_a(FP16MAC4_io_a),
    .io_b(FP16MAC4_io_b),
    .io_c(FP16MAC4_io_c),
    .io_out(FP16MAC4_io_out)
  );
  tanh_Unit tanh ( // @[Unit.scala 527:20]
    .io_input(tanh_io_input),
    .io_output(tanh_io_output)
  );
  assign io_output = reg_output; // @[Unit.scala 550:15]
  assign FP16MAC1_io_a = io_Rt_input; // @[Unit.scala 520:17]
  assign FP16MAC1_io_b = io_Uhht_1_input; // @[Unit.scala 521:17]
  assign FP16MAC1_io_c = io_Whxt_input; // @[Unit.scala 522:17]
  assign FP16MAC2_io_a = {reg_Zt_inv_hi,reg_Zt_inv_lo}; // @[Cat.scala 30:58]
  assign FP16MAC2_io_b = 16'h3c00; // @[Unit.scala 534:17]
  assign FP16MAC2_io_c = 16'h3c00; // @[Unit.scala 535:17]
  assign FP16MAC3_io_a = reg_Zt; // @[Unit.scala 539:17]
  assign FP16MAC3_io_b = reg_ht_1; // @[Unit.scala 540:17]
  assign FP16MAC3_io_c = 16'h0; // @[Unit.scala 541:17]
  assign FP16MAC4_io_a = reg_tanh; // @[Unit.scala 545:17]
  assign FP16MAC4_io_b = reg_1_Zt; // @[Unit.scala 546:17]
  assign FP16MAC4_io_c = reg_Zt_ht_1; // @[Unit.scala 547:17]
  assign tanh_io_input = reg_before_tanh; // @[Unit.scala 528:17]
  always @(posedge clock) begin
    if (reset) begin // @[Unit.scala 493:32]
      reg_before_tanh <= 16'h0; // @[Unit.scala 493:32]
    end else begin
      reg_before_tanh <= FP16MAC1_io_out; // @[Unit.scala 523:19]
    end
    if (reset) begin // @[Unit.scala 494:30]
      reg_Zt <= 16'h0; // @[Unit.scala 494:30]
    end else begin
      reg_Zt <= io_Zt_input; // @[Unit.scala 525:17]
    end
    if (reset) begin // @[Unit.scala 495:30]
      reg_ht_1 <= 16'h0; // @[Unit.scala 495:30]
    end else begin
      reg_ht_1 <= io_ht_1_input; // @[Unit.scala 526:17]
    end
    if (reset) begin // @[Unit.scala 496:30]
      reg_tanh <= 16'h0; // @[Unit.scala 496:30]
    end else begin
      reg_tanh <= tanh_io_output; // @[Unit.scala 529:17]
    end
    if (reset) begin // @[Unit.scala 497:30]
      reg_1_Zt <= 16'h0; // @[Unit.scala 497:30]
    end else begin
      reg_1_Zt <= FP16MAC2_io_out; // @[Unit.scala 536:17]
    end
    if (reset) begin // @[Unit.scala 498:30]
      reg_Zt_ht_1 <= 16'h0; // @[Unit.scala 498:30]
    end else begin
      reg_Zt_ht_1 <= FP16MAC3_io_out; // @[Unit.scala 542:17]
    end
    if (reset) begin // @[Unit.scala 499:30]
      reg_output <= 16'h0; // @[Unit.scala 499:30]
    end else begin
      reg_output <= FP16MAC4_io_out; // @[Unit.scala 548:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_before_tanh = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  reg_Zt = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  reg_ht_1 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  reg_tanh = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  reg_1_Zt = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  reg_Zt_ht_1 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  reg_output = _RAND_6[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module accumulator_registers_4(
  input         clock,
  input         reset,
  output [15:0] io_rdData,
  input         io_wrEna,
  input  [15:0] io_wrData,
  input  [3:0]  io_wrAddr
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] FP16MAC_io_a; // @[Unit.scala 389:23]
  wire [15:0] FP16MAC_io_b; // @[Unit.scala 389:23]
  wire [15:0] FP16MAC_io_c; // @[Unit.scala 389:23]
  wire [15:0] FP16MAC_io_out; // @[Unit.scala 389:23]
  reg [15:0] register_0; // @[Unit.scala 386:25]
  reg [15:0] register_1; // @[Unit.scala 386:25]
  reg [15:0] register_2; // @[Unit.scala 386:25]
  reg [15:0] register_3; // @[Unit.scala 386:25]
  reg [15:0] register_4; // @[Unit.scala 386:25]
  reg [15:0] register_5; // @[Unit.scala 386:25]
  wire [15:0] _GEN_7 = 3'h1 == io_wrAddr[2:0] ? register_1 : register_0; // @[Unit.scala 398:18 Unit.scala 398:18]
  wire [15:0] _GEN_8 = 3'h2 == io_wrAddr[2:0] ? register_2 : _GEN_7; // @[Unit.scala 398:18 Unit.scala 398:18]
  wire [15:0] _GEN_9 = 3'h3 == io_wrAddr[2:0] ? register_3 : _GEN_8; // @[Unit.scala 398:18 Unit.scala 398:18]
  wire [15:0] _GEN_10 = 3'h4 == io_wrAddr[2:0] ? register_4 : _GEN_9; // @[Unit.scala 398:18 Unit.scala 398:18]
  wire [15:0] _GEN_11 = 3'h5 == io_wrAddr[2:0] ? register_5 : _GEN_10; // @[Unit.scala 398:18 Unit.scala 398:18]
  wire [15:0] _register_T = FP16MAC_io_out; // @[Unit.scala 399:25 Unit.scala 399:25]
  wire [13:0] _GEN_19 = io_wrEna ? 14'h3c00 : 14'h0; // @[Unit.scala 395:17 Unit.scala 397:18 Unit.scala 403:20]
  FP16MulAdder FP16MAC ( // @[Unit.scala 389:23]
    .io_a(FP16MAC_io_a),
    .io_b(FP16MAC_io_b),
    .io_c(FP16MAC_io_c),
    .io_out(FP16MAC_io_out)
  );
  assign io_rdData = register_0; // @[Unit.scala 394:13 Unit.scala 394:13]
  assign FP16MAC_io_a = io_wrEna ? io_wrData : 16'h0; // @[Unit.scala 395:17 Unit.scala 396:18 Unit.scala 402:20]
  assign FP16MAC_io_b = {{2'd0}, _GEN_19}; // @[Unit.scala 395:17 Unit.scala 397:18 Unit.scala 403:20]
  assign FP16MAC_io_c = io_wrEna ? _GEN_11 : 16'h0; // @[Unit.scala 395:17 Unit.scala 398:18 Unit.scala 404:20]
  always @(posedge clock) begin
    if (reset) begin // @[Unit.scala 386:25]
      register_0 <= 16'h0; // @[Unit.scala 386:25]
    end else if (io_wrEna) begin // @[Unit.scala 395:17]
      if (3'h0 == io_wrAddr[2:0]) begin // @[Unit.scala 399:25]
        register_0 <= _register_T; // @[Unit.scala 399:25]
      end
    end
    if (reset) begin // @[Unit.scala 386:25]
      register_1 <= 16'h0; // @[Unit.scala 386:25]
    end else if (io_wrEna) begin // @[Unit.scala 395:17]
      if (3'h1 == io_wrAddr[2:0]) begin // @[Unit.scala 399:25]
        register_1 <= _register_T; // @[Unit.scala 399:25]
      end
    end
    if (reset) begin // @[Unit.scala 386:25]
      register_2 <= 16'h0; // @[Unit.scala 386:25]
    end else if (io_wrEna) begin // @[Unit.scala 395:17]
      if (3'h2 == io_wrAddr[2:0]) begin // @[Unit.scala 399:25]
        register_2 <= _register_T; // @[Unit.scala 399:25]
      end
    end
    if (reset) begin // @[Unit.scala 386:25]
      register_3 <= 16'h0; // @[Unit.scala 386:25]
    end else if (io_wrEna) begin // @[Unit.scala 395:17]
      if (3'h3 == io_wrAddr[2:0]) begin // @[Unit.scala 399:25]
        register_3 <= _register_T; // @[Unit.scala 399:25]
      end
    end
    if (reset) begin // @[Unit.scala 386:25]
      register_4 <= 16'h0; // @[Unit.scala 386:25]
    end else if (io_wrEna) begin // @[Unit.scala 395:17]
      if (3'h4 == io_wrAddr[2:0]) begin // @[Unit.scala 399:25]
        register_4 <= _register_T; // @[Unit.scala 399:25]
      end
    end
    if (reset) begin // @[Unit.scala 386:25]
      register_5 <= 16'h0; // @[Unit.scala 386:25]
    end else if (io_wrEna) begin // @[Unit.scala 395:17]
      if (3'h5 == io_wrAddr[2:0]) begin // @[Unit.scala 399:25]
        register_5 <= _register_T; // @[Unit.scala 399:25]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  register_0 = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  register_1 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  register_2 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  register_3 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  register_4 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  register_5 = _RAND_5[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Top(
  input         clock,
  input         reset,
  input         io_Start,
  input  [15:0] io_Input_Data,
  input         io_Input_Valid,
  output        io_Input_Ready,
  output [15:0] io_Output_Data,
  input         io_Output_Ready
);
  wire  L1_Memory_top_0_clock; // @[Top.scala 17:42]
  wire [11:0] L1_Memory_top_0_io_rdAddr; // @[Top.scala 17:42]
  wire [15:0] L1_Memory_top_0_io_rdData; // @[Top.scala 17:42]
  wire  L1_Memory_top_0_io_wrEna; // @[Top.scala 17:42]
  wire [15:0] L1_Memory_top_0_io_wrData; // @[Top.scala 17:42]
  wire [11:0] L1_Memory_top_0_io_wrAddr; // @[Top.scala 17:42]
  wire  L1_Memory_top_1_clock; // @[Top.scala 17:42]
  wire [11:0] L1_Memory_top_1_io_rdAddr; // @[Top.scala 17:42]
  wire [15:0] L1_Memory_top_1_io_rdData; // @[Top.scala 17:42]
  wire  L1_Memory_top_1_io_wrEna; // @[Top.scala 17:42]
  wire [15:0] L1_Memory_top_1_io_wrData; // @[Top.scala 17:42]
  wire [11:0] L1_Memory_top_1_io_wrAddr; // @[Top.scala 17:42]
  wire  L1_Memory_top_2_clock; // @[Top.scala 17:42]
  wire [11:0] L1_Memory_top_2_io_rdAddr; // @[Top.scala 17:42]
  wire [15:0] L1_Memory_top_2_io_rdData; // @[Top.scala 17:42]
  wire  L1_Memory_top_2_io_wrEna; // @[Top.scala 17:42]
  wire [15:0] L1_Memory_top_2_io_wrData; // @[Top.scala 17:42]
  wire [11:0] L1_Memory_top_2_io_wrAddr; // @[Top.scala 17:42]
  wire  L1_Memory_top_3_clock; // @[Top.scala 17:42]
  wire [11:0] L1_Memory_top_3_io_rdAddr; // @[Top.scala 17:42]
  wire [15:0] L1_Memory_top_3_io_rdData; // @[Top.scala 17:42]
  wire  L1_Memory_top_3_io_wrEna; // @[Top.scala 17:42]
  wire [15:0] L1_Memory_top_3_io_wrData; // @[Top.scala 17:42]
  wire [11:0] L1_Memory_top_3_io_wrAddr; // @[Top.scala 17:42]
  wire  L1_Memory_top_4_clock; // @[Top.scala 17:42]
  wire [11:0] L1_Memory_top_4_io_rdAddr; // @[Top.scala 17:42]
  wire [15:0] L1_Memory_top_4_io_rdData; // @[Top.scala 17:42]
  wire  L1_Memory_top_4_io_wrEna; // @[Top.scala 17:42]
  wire [15:0] L1_Memory_top_4_io_wrData; // @[Top.scala 17:42]
  wire [11:0] L1_Memory_top_4_io_wrAddr; // @[Top.scala 17:42]
  wire  L1_Memory_top_5_clock; // @[Top.scala 17:42]
  wire [11:0] L1_Memory_top_5_io_rdAddr; // @[Top.scala 17:42]
  wire [15:0] L1_Memory_top_5_io_rdData; // @[Top.scala 17:42]
  wire  L1_Memory_top_5_io_wrEna; // @[Top.scala 17:42]
  wire [15:0] L1_Memory_top_5_io_wrData; // @[Top.scala 17:42]
  wire [11:0] L1_Memory_top_5_io_wrAddr; // @[Top.scala 17:42]
  wire  L1_Memory_top_6_clock; // @[Top.scala 17:42]
  wire [11:0] L1_Memory_top_6_io_rdAddr; // @[Top.scala 17:42]
  wire [15:0] L1_Memory_top_6_io_rdData; // @[Top.scala 17:42]
  wire  L1_Memory_top_6_io_wrEna; // @[Top.scala 17:42]
  wire [15:0] L1_Memory_top_6_io_wrData; // @[Top.scala 17:42]
  wire [11:0] L1_Memory_top_6_io_wrAddr; // @[Top.scala 17:42]
  wire  L1_Memory_top_7_clock; // @[Top.scala 17:42]
  wire [11:0] L1_Memory_top_7_io_rdAddr; // @[Top.scala 17:42]
  wire [15:0] L1_Memory_top_7_io_rdData; // @[Top.scala 17:42]
  wire  L1_Memory_top_7_io_wrEna; // @[Top.scala 17:42]
  wire [15:0] L1_Memory_top_7_io_wrData; // @[Top.scala 17:42]
  wire [11:0] L1_Memory_top_7_io_wrAddr; // @[Top.scala 17:42]
  wire  L1_Memory_top_8_clock; // @[Top.scala 17:42]
  wire [11:0] L1_Memory_top_8_io_rdAddr; // @[Top.scala 17:42]
  wire [15:0] L1_Memory_top_8_io_rdData; // @[Top.scala 17:42]
  wire  L1_Memory_top_8_io_wrEna; // @[Top.scala 17:42]
  wire [15:0] L1_Memory_top_8_io_wrData; // @[Top.scala 17:42]
  wire [11:0] L1_Memory_top_8_io_wrAddr; // @[Top.scala 17:42]
  wire  L1_Memory_top_9_clock; // @[Top.scala 17:42]
  wire [11:0] L1_Memory_top_9_io_rdAddr; // @[Top.scala 17:42]
  wire [15:0] L1_Memory_top_9_io_rdData; // @[Top.scala 17:42]
  wire  L1_Memory_top_9_io_wrEna; // @[Top.scala 17:42]
  wire [15:0] L1_Memory_top_9_io_wrData; // @[Top.scala 17:42]
  wire [11:0] L1_Memory_top_9_io_wrAddr; // @[Top.scala 17:42]
  wire  L1_Memory_top_10_clock; // @[Top.scala 17:42]
  wire [11:0] L1_Memory_top_10_io_rdAddr; // @[Top.scala 17:42]
  wire [15:0] L1_Memory_top_10_io_rdData; // @[Top.scala 17:42]
  wire  L1_Memory_top_10_io_wrEna; // @[Top.scala 17:42]
  wire [15:0] L1_Memory_top_10_io_wrData; // @[Top.scala 17:42]
  wire [11:0] L1_Memory_top_10_io_wrAddr; // @[Top.scala 17:42]
  wire  L1_Memory_top_11_clock; // @[Top.scala 17:42]
  wire [11:0] L1_Memory_top_11_io_rdAddr; // @[Top.scala 17:42]
  wire [15:0] L1_Memory_top_11_io_rdData; // @[Top.scala 17:42]
  wire  L1_Memory_top_11_io_wrEna; // @[Top.scala 17:42]
  wire [15:0] L1_Memory_top_11_io_wrData; // @[Top.scala 17:42]
  wire [11:0] L1_Memory_top_11_io_wrAddr; // @[Top.scala 17:42]
  wire  PEArray_top_clock; // @[Top.scala 18:27]
  wire  PEArray_top_reset; // @[Top.scala 18:27]
  wire [15:0] PEArray_top_io_From_above_0; // @[Top.scala 18:27]
  wire [15:0] PEArray_top_io_From_above_1; // @[Top.scala 18:27]
  wire [15:0] PEArray_top_io_From_above_2; // @[Top.scala 18:27]
  wire [15:0] PEArray_top_io_From_above_3; // @[Top.scala 18:27]
  wire [15:0] PEArray_top_io_From_above_4; // @[Top.scala 18:27]
  wire [15:0] PEArray_top_io_From_above_5; // @[Top.scala 18:27]
  wire [15:0] PEArray_top_io_From_above_6; // @[Top.scala 18:27]
  wire [15:0] PEArray_top_io_From_above_7; // @[Top.scala 18:27]
  wire [15:0] PEArray_top_io_From_above_8; // @[Top.scala 18:27]
  wire [15:0] PEArray_top_io_From_above_9; // @[Top.scala 18:27]
  wire [15:0] PEArray_top_io_From_above_10; // @[Top.scala 18:27]
  wire [15:0] PEArray_top_io_From_above_11; // @[Top.scala 18:27]
  wire [11:0] PEArray_top_io_PE_control_0_mask; // @[Top.scala 18:27]
  wire [11:0] PEArray_top_io_PE_control_1_mask; // @[Top.scala 18:27]
  wire [2:0] PEArray_top_io_PE_control_2_control; // @[Top.scala 18:27]
  wire [9:0] PEArray_top_io_PE_control_2_count; // @[Top.scala 18:27]
  wire [5:0] PEArray_top_io_PE_control_2_L0index; // @[Top.scala 18:27]
  wire [11:0] PEArray_top_io_PE_control_2_mask; // @[Top.scala 18:27]
  wire [7:0] PEArray_top_io_PE_control_2_gru_out_width; // @[Top.scala 18:27]
  wire [3:0] PEArray_top_io_rd_data_mux; // @[Top.scala 18:27]
  wire [15:0] PEArray_top_io_To_below_0; // @[Top.scala 18:27]
  wire [15:0] PEArray_top_io_To_below_1; // @[Top.scala 18:27]
  wire [15:0] PEArray_top_io_To_below_2; // @[Top.scala 18:27]
  wire [15:0] PEArray_top_io_To_below_3; // @[Top.scala 18:27]
  wire [15:0] PEArray_top_io_To_below_4; // @[Top.scala 18:27]
  wire [15:0] PEArray_top_io_To_below_5; // @[Top.scala 18:27]
  wire [15:0] PEArray_top_io_To_below_6; // @[Top.scala 18:27]
  wire [15:0] PEArray_top_io_To_below_7; // @[Top.scala 18:27]
  wire [15:0] PEArray_top_io_To_below_8; // @[Top.scala 18:27]
  wire [15:0] PEArray_top_io_To_below_9; // @[Top.scala 18:27]
  wire [15:0] PEArray_top_io_To_below_10; // @[Top.scala 18:27]
  wire [15:0] PEArray_top_io_To_below_11; // @[Top.scala 18:27]
  wire [15:0] PEArray_top_io_To_right_2; // @[Top.scala 18:27]
  wire  FSM_top_clock; // @[Top.scala 19:23]
  wire  FSM_top_reset; // @[Top.scala 19:23]
  wire  FSM_top_io_Start; // @[Top.scala 19:23]
  wire [15:0] FSM_top_io_Input_Data; // @[Top.scala 19:23]
  wire  FSM_top_io_Input_Valid; // @[Top.scala 19:23]
  wire  FSM_top_io_Input_Ready; // @[Top.scala 19:23]
  wire [15:0] FSM_top_io_L1_wr_data; // @[Top.scala 19:23]
  wire  FSM_top_io_To_L1_control; // @[Top.scala 19:23]
  wire [11:0] FSM_top_io_L1_rd_addr_0; // @[Top.scala 19:23]
  wire [11:0] FSM_top_io_L1_rd_addr_1; // @[Top.scala 19:23]
  wire [11:0] FSM_top_io_L1_rd_addr_2; // @[Top.scala 19:23]
  wire [11:0] FSM_top_io_L1_rd_addr_3; // @[Top.scala 19:23]
  wire [11:0] FSM_top_io_L1_rd_addr_4; // @[Top.scala 19:23]
  wire [11:0] FSM_top_io_L1_rd_addr_5; // @[Top.scala 19:23]
  wire [11:0] FSM_top_io_L1_rd_addr_6; // @[Top.scala 19:23]
  wire [11:0] FSM_top_io_L1_rd_addr_7; // @[Top.scala 19:23]
  wire [11:0] FSM_top_io_L1_rd_addr_8; // @[Top.scala 19:23]
  wire [11:0] FSM_top_io_L1_rd_addr_9; // @[Top.scala 19:23]
  wire [11:0] FSM_top_io_L1_rd_addr_10; // @[Top.scala 19:23]
  wire [11:0] FSM_top_io_L1_rd_addr_11; // @[Top.scala 19:23]
  wire [3:0] FSM_top_io_PE_rd_data_mux; // @[Top.scala 19:23]
  wire [11:0] FSM_top_io_L1_wr_addr_0; // @[Top.scala 19:23]
  wire [11:0] FSM_top_io_L1_wr_addr_1; // @[Top.scala 19:23]
  wire [11:0] FSM_top_io_L1_wr_addr_2; // @[Top.scala 19:23]
  wire [11:0] FSM_top_io_L1_wr_addr_3; // @[Top.scala 19:23]
  wire [11:0] FSM_top_io_L1_wr_addr_4; // @[Top.scala 19:23]
  wire [11:0] FSM_top_io_L1_wr_addr_5; // @[Top.scala 19:23]
  wire [11:0] FSM_top_io_L1_wr_addr_6; // @[Top.scala 19:23]
  wire [11:0] FSM_top_io_L1_wr_addr_7; // @[Top.scala 19:23]
  wire [11:0] FSM_top_io_L1_wr_addr_8; // @[Top.scala 19:23]
  wire [11:0] FSM_top_io_L1_wr_addr_9; // @[Top.scala 19:23]
  wire [11:0] FSM_top_io_L1_wr_addr_10; // @[Top.scala 19:23]
  wire [11:0] FSM_top_io_L1_wr_addr_11; // @[Top.scala 19:23]
  wire  FSM_top_io_L1_wrEna_0; // @[Top.scala 19:23]
  wire  FSM_top_io_L1_wrEna_1; // @[Top.scala 19:23]
  wire  FSM_top_io_L1_wrEna_2; // @[Top.scala 19:23]
  wire  FSM_top_io_L1_wrEna_3; // @[Top.scala 19:23]
  wire  FSM_top_io_L1_wrEna_4; // @[Top.scala 19:23]
  wire  FSM_top_io_L1_wrEna_5; // @[Top.scala 19:23]
  wire  FSM_top_io_L1_wrEna_6; // @[Top.scala 19:23]
  wire  FSM_top_io_L1_wrEna_7; // @[Top.scala 19:23]
  wire  FSM_top_io_L1_wrEna_8; // @[Top.scala 19:23]
  wire  FSM_top_io_L1_wrEna_9; // @[Top.scala 19:23]
  wire  FSM_top_io_L1_wrEna_10; // @[Top.scala 19:23]
  wire  FSM_top_io_L1_wrEna_11; // @[Top.scala 19:23]
  wire [11:0] FSM_top_io_PEArray_ctrl_0_mask; // @[Top.scala 19:23]
  wire [11:0] FSM_top_io_PEArray_ctrl_1_mask; // @[Top.scala 19:23]
  wire [2:0] FSM_top_io_PEArray_ctrl_2_control; // @[Top.scala 19:23]
  wire [9:0] FSM_top_io_PEArray_ctrl_2_count; // @[Top.scala 19:23]
  wire [5:0] FSM_top_io_PEArray_ctrl_2_L0index; // @[Top.scala 19:23]
  wire [11:0] FSM_top_io_PEArray_ctrl_2_mask; // @[Top.scala 19:23]
  wire [7:0] FSM_top_io_PEArray_ctrl_2_gru_out_width; // @[Top.scala 19:23]
  wire [1:0] FSM_top_io_BNArray_ctrl_0; // @[Top.scala 19:23]
  wire [1:0] FSM_top_io_BNArray_ctrl_1; // @[Top.scala 19:23]
  wire [1:0] FSM_top_io_BNArray_ctrl_2; // @[Top.scala 19:23]
  wire [1:0] FSM_top_io_BNArray_ctrl_3; // @[Top.scala 19:23]
  wire [1:0] FSM_top_io_BNArray_ctrl_4; // @[Top.scala 19:23]
  wire [1:0] FSM_top_io_BNArray_ctrl_5; // @[Top.scala 19:23]
  wire [1:0] FSM_top_io_BNArray_ctrl_6; // @[Top.scala 19:23]
  wire [1:0] FSM_top_io_BNArray_ctrl_7; // @[Top.scala 19:23]
  wire [1:0] FSM_top_io_BNArray_ctrl_8; // @[Top.scala 19:23]
  wire [1:0] FSM_top_io_BNArray_ctrl_9; // @[Top.scala 19:23]
  wire [1:0] FSM_top_io_BNArray_ctrl_10; // @[Top.scala 19:23]
  wire [1:0] FSM_top_io_BNArray_ctrl_11; // @[Top.scala 19:23]
  wire [1:0] FSM_top_io_BN_Unit_ctrl; // @[Top.scala 19:23]
  wire  FSM_top_io_Relu6Array_ctrl_0; // @[Top.scala 19:23]
  wire  FSM_top_io_Relu6Array_ctrl_1; // @[Top.scala 19:23]
  wire  FSM_top_io_Relu6Array_ctrl_2; // @[Top.scala 19:23]
  wire  FSM_top_io_Relu6Array_ctrl_3; // @[Top.scala 19:23]
  wire  FSM_top_io_Relu6Array_ctrl_4; // @[Top.scala 19:23]
  wire  FSM_top_io_Relu6Array_ctrl_5; // @[Top.scala 19:23]
  wire  FSM_top_io_Relu6Array_ctrl_6; // @[Top.scala 19:23]
  wire  FSM_top_io_Relu6Array_ctrl_7; // @[Top.scala 19:23]
  wire  FSM_top_io_Relu6Array_ctrl_8; // @[Top.scala 19:23]
  wire  FSM_top_io_Relu6Array_ctrl_9; // @[Top.scala 19:23]
  wire  FSM_top_io_Relu6Array_ctrl_10; // @[Top.scala 19:23]
  wire  FSM_top_io_Relu6Array_ctrl_11; // @[Top.scala 19:23]
  wire [1:0] FSM_top_io_PE_above_data_ctrl; // @[Top.scala 19:23]
  wire [1:0] FSM_top_io_Activation_ctrl; // @[Top.scala 19:23]
  wire [2:0] FSM_top_io_Ht_to_PE_control; // @[Top.scala 19:23]
  wire  FSM_top_io_Ht_wrEna; // @[Top.scala 19:23]
  wire [5:0] FSM_top_io_Ht_wrAddr; // @[Top.scala 19:23]
  wire [5:0] FSM_top_io_Zt_rdAddr; // @[Top.scala 19:23]
  wire  FSM_top_io_Zt_wrEna; // @[Top.scala 19:23]
  wire [5:0] FSM_top_io_Zt_wrAddr; // @[Top.scala 19:23]
  wire [5:0] FSM_top_io_Rt_rdAddr; // @[Top.scala 19:23]
  wire  FSM_top_io_Rt_wrEna; // @[Top.scala 19:23]
  wire [5:0] FSM_top_io_Rt_wrAddr; // @[Top.scala 19:23]
  wire [5:0] FSM_top_io_WhXt_rdAddr; // @[Top.scala 19:23]
  wire  FSM_top_io_WhXt_wrEna; // @[Top.scala 19:23]
  wire [5:0] FSM_top_io_WhXt_wrAddr; // @[Top.scala 19:23]
  wire [5:0] FSM_top_io_Uhht_1_rdAddr; // @[Top.scala 19:23]
  wire  FSM_top_io_Uhht_1_wrEna; // @[Top.scala 19:23]
  wire [5:0] FSM_top_io_Uhht_1_wrAddr; // @[Top.scala 19:23]
  wire [2:0] FSM_top_io_FC_temp_to_PE_control; // @[Top.scala 19:23]
  wire  FSM_top_io_FC_temp_wrEna; // @[Top.scala 19:23]
  wire [5:0] FSM_top_io_FC_temp_wrAddr; // @[Top.scala 19:23]
  wire  FSM_top_io_Result_wrEna; // @[Top.scala 19:23]
  wire [3:0] FSM_top_io_Result_wrAddr; // @[Top.scala 19:23]
  wire  BN_Array_below_clock; // @[Top.scala 21:30]
  wire  BN_Array_below_reset; // @[Top.scala 21:30]
  wire [15:0] BN_Array_below_io_from_PE_0; // @[Top.scala 21:30]
  wire [15:0] BN_Array_below_io_from_PE_1; // @[Top.scala 21:30]
  wire [15:0] BN_Array_below_io_from_PE_2; // @[Top.scala 21:30]
  wire [15:0] BN_Array_below_io_from_PE_3; // @[Top.scala 21:30]
  wire [15:0] BN_Array_below_io_from_PE_4; // @[Top.scala 21:30]
  wire [15:0] BN_Array_below_io_from_PE_5; // @[Top.scala 21:30]
  wire [15:0] BN_Array_below_io_from_PE_6; // @[Top.scala 21:30]
  wire [15:0] BN_Array_below_io_from_PE_7; // @[Top.scala 21:30]
  wire [15:0] BN_Array_below_io_from_PE_8; // @[Top.scala 21:30]
  wire [15:0] BN_Array_below_io_from_PE_9; // @[Top.scala 21:30]
  wire [15:0] BN_Array_below_io_from_PE_10; // @[Top.scala 21:30]
  wire [15:0] BN_Array_below_io_from_PE_11; // @[Top.scala 21:30]
  wire [1:0] BN_Array_below_io_control_0; // @[Top.scala 21:30]
  wire [1:0] BN_Array_below_io_control_1; // @[Top.scala 21:30]
  wire [1:0] BN_Array_below_io_control_2; // @[Top.scala 21:30]
  wire [1:0] BN_Array_below_io_control_3; // @[Top.scala 21:30]
  wire [1:0] BN_Array_below_io_control_4; // @[Top.scala 21:30]
  wire [1:0] BN_Array_below_io_control_5; // @[Top.scala 21:30]
  wire [1:0] BN_Array_below_io_control_6; // @[Top.scala 21:30]
  wire [1:0] BN_Array_below_io_control_7; // @[Top.scala 21:30]
  wire [1:0] BN_Array_below_io_control_8; // @[Top.scala 21:30]
  wire [1:0] BN_Array_below_io_control_9; // @[Top.scala 21:30]
  wire [1:0] BN_Array_below_io_control_10; // @[Top.scala 21:30]
  wire [1:0] BN_Array_below_io_control_11; // @[Top.scala 21:30]
  wire [15:0] BN_Array_below_io_to_Relu6_0; // @[Top.scala 21:30]
  wire [15:0] BN_Array_below_io_to_Relu6_1; // @[Top.scala 21:30]
  wire [15:0] BN_Array_below_io_to_Relu6_2; // @[Top.scala 21:30]
  wire [15:0] BN_Array_below_io_to_Relu6_3; // @[Top.scala 21:30]
  wire [15:0] BN_Array_below_io_to_Relu6_4; // @[Top.scala 21:30]
  wire [15:0] BN_Array_below_io_to_Relu6_5; // @[Top.scala 21:30]
  wire [15:0] BN_Array_below_io_to_Relu6_6; // @[Top.scala 21:30]
  wire [15:0] BN_Array_below_io_to_Relu6_7; // @[Top.scala 21:30]
  wire [15:0] BN_Array_below_io_to_Relu6_8; // @[Top.scala 21:30]
  wire [15:0] BN_Array_below_io_to_Relu6_9; // @[Top.scala 21:30]
  wire [15:0] BN_Array_below_io_to_Relu6_10; // @[Top.scala 21:30]
  wire [15:0] BN_Array_below_io_to_Relu6_11; // @[Top.scala 21:30]
  wire [15:0] Relu6_Array_io_input_0; // @[Top.scala 22:27]
  wire [15:0] Relu6_Array_io_input_1; // @[Top.scala 22:27]
  wire [15:0] Relu6_Array_io_input_2; // @[Top.scala 22:27]
  wire [15:0] Relu6_Array_io_input_3; // @[Top.scala 22:27]
  wire [15:0] Relu6_Array_io_input_4; // @[Top.scala 22:27]
  wire [15:0] Relu6_Array_io_input_5; // @[Top.scala 22:27]
  wire [15:0] Relu6_Array_io_input_6; // @[Top.scala 22:27]
  wire [15:0] Relu6_Array_io_input_7; // @[Top.scala 22:27]
  wire [15:0] Relu6_Array_io_input_8; // @[Top.scala 22:27]
  wire [15:0] Relu6_Array_io_input_9; // @[Top.scala 22:27]
  wire [15:0] Relu6_Array_io_input_10; // @[Top.scala 22:27]
  wire [15:0] Relu6_Array_io_input_11; // @[Top.scala 22:27]
  wire  Relu6_Array_io_control_0; // @[Top.scala 22:27]
  wire  Relu6_Array_io_control_1; // @[Top.scala 22:27]
  wire  Relu6_Array_io_control_2; // @[Top.scala 22:27]
  wire  Relu6_Array_io_control_3; // @[Top.scala 22:27]
  wire  Relu6_Array_io_control_4; // @[Top.scala 22:27]
  wire  Relu6_Array_io_control_5; // @[Top.scala 22:27]
  wire  Relu6_Array_io_control_6; // @[Top.scala 22:27]
  wire  Relu6_Array_io_control_7; // @[Top.scala 22:27]
  wire  Relu6_Array_io_control_8; // @[Top.scala 22:27]
  wire  Relu6_Array_io_control_9; // @[Top.scala 22:27]
  wire  Relu6_Array_io_control_10; // @[Top.scala 22:27]
  wire  Relu6_Array_io_control_11; // @[Top.scala 22:27]
  wire [15:0] Relu6_Array_io_output_0; // @[Top.scala 22:27]
  wire [15:0] Relu6_Array_io_output_1; // @[Top.scala 22:27]
  wire [15:0] Relu6_Array_io_output_2; // @[Top.scala 22:27]
  wire [15:0] Relu6_Array_io_output_3; // @[Top.scala 22:27]
  wire [15:0] Relu6_Array_io_output_4; // @[Top.scala 22:27]
  wire [15:0] Relu6_Array_io_output_5; // @[Top.scala 22:27]
  wire [15:0] Relu6_Array_io_output_6; // @[Top.scala 22:27]
  wire [15:0] Relu6_Array_io_output_7; // @[Top.scala 22:27]
  wire [15:0] Relu6_Array_io_output_8; // @[Top.scala 22:27]
  wire [15:0] Relu6_Array_io_output_9; // @[Top.scala 22:27]
  wire [15:0] Relu6_Array_io_output_10; // @[Top.scala 22:27]
  wire [15:0] Relu6_Array_io_output_11; // @[Top.scala 22:27]
  wire  BNUnit_right_clock; // @[Top.scala 23:28]
  wire  BNUnit_right_reset; // @[Top.scala 23:28]
  wire [15:0] BNUnit_right_io_input; // @[Top.scala 23:28]
  wire [1:0] BNUnit_right_io_control; // @[Top.scala 23:28]
  wire [15:0] BNUnit_right_io_output; // @[Top.scala 23:28]
  wire  Activation_clock; // @[Top.scala 24:26]
  wire  Activation_reset; // @[Top.scala 24:26]
  wire [15:0] Activation_io_input; // @[Top.scala 24:26]
  wire [1:0] Activation_io_control; // @[Top.scala 24:26]
  wire [15:0] Activation_io_output; // @[Top.scala 24:26]
  wire  Zt_clock; // @[Top.scala 26:18]
  wire  Zt_reset; // @[Top.scala 26:18]
  wire [5:0] Zt_io_rdAddr; // @[Top.scala 26:18]
  wire [15:0] Zt_io_rdData; // @[Top.scala 26:18]
  wire  Zt_io_wrEna; // @[Top.scala 26:18]
  wire [15:0] Zt_io_wrData; // @[Top.scala 26:18]
  wire [5:0] Zt_io_wrAddr; // @[Top.scala 26:18]
  wire  Rt_clock; // @[Top.scala 27:18]
  wire  Rt_reset; // @[Top.scala 27:18]
  wire [5:0] Rt_io_rdAddr; // @[Top.scala 27:18]
  wire [15:0] Rt_io_rdData; // @[Top.scala 27:18]
  wire  Rt_io_wrEna; // @[Top.scala 27:18]
  wire [15:0] Rt_io_wrData; // @[Top.scala 27:18]
  wire [5:0] Rt_io_wrAddr; // @[Top.scala 27:18]
  wire  WhXt_clock; // @[Top.scala 28:20]
  wire  WhXt_reset; // @[Top.scala 28:20]
  wire [5:0] WhXt_io_rdAddr; // @[Top.scala 28:20]
  wire [15:0] WhXt_io_rdData; // @[Top.scala 28:20]
  wire  WhXt_io_wrEna; // @[Top.scala 28:20]
  wire [15:0] WhXt_io_wrData; // @[Top.scala 28:20]
  wire [5:0] WhXt_io_wrAddr; // @[Top.scala 28:20]
  wire  Uhht_1_clock; // @[Top.scala 29:22]
  wire  Uhht_1_reset; // @[Top.scala 29:22]
  wire [5:0] Uhht_1_io_rdAddr; // @[Top.scala 29:22]
  wire [15:0] Uhht_1_io_rdData; // @[Top.scala 29:22]
  wire  Uhht_1_io_wrEna; // @[Top.scala 29:22]
  wire [15:0] Uhht_1_io_wrData; // @[Top.scala 29:22]
  wire [5:0] Uhht_1_io_wrAddr; // @[Top.scala 29:22]
  wire  Ht_clock; // @[Top.scala 30:18]
  wire  Ht_reset; // @[Top.scala 30:18]
  wire [15:0] Ht_io_to_PE_0; // @[Top.scala 30:18]
  wire [15:0] Ht_io_to_PE_1; // @[Top.scala 30:18]
  wire [15:0] Ht_io_to_PE_2; // @[Top.scala 30:18]
  wire [15:0] Ht_io_to_PE_3; // @[Top.scala 30:18]
  wire [15:0] Ht_io_to_PE_4; // @[Top.scala 30:18]
  wire [15:0] Ht_io_to_PE_5; // @[Top.scala 30:18]
  wire [15:0] Ht_io_to_PE_6; // @[Top.scala 30:18]
  wire [15:0] Ht_io_to_PE_7; // @[Top.scala 30:18]
  wire [15:0] Ht_io_to_PE_8; // @[Top.scala 30:18]
  wire [15:0] Ht_io_to_PE_9; // @[Top.scala 30:18]
  wire [15:0] Ht_io_to_PE_10; // @[Top.scala 30:18]
  wire [15:0] Ht_io_to_PE_11; // @[Top.scala 30:18]
  wire [2:0] Ht_io_to_PE_control; // @[Top.scala 30:18]
  wire [15:0] Ht_io_rdData; // @[Top.scala 30:18]
  wire  Ht_io_wrEna; // @[Top.scala 30:18]
  wire [15:0] Ht_io_wrData; // @[Top.scala 30:18]
  wire [5:0] Ht_io_wrAddr; // @[Top.scala 30:18]
  wire  EW_clock; // @[Top.scala 31:18]
  wire  EW_reset; // @[Top.scala 31:18]
  wire [15:0] EW_io_ht_1_input; // @[Top.scala 31:18]
  wire [15:0] EW_io_Zt_input; // @[Top.scala 31:18]
  wire [15:0] EW_io_Rt_input; // @[Top.scala 31:18]
  wire [15:0] EW_io_Whxt_input; // @[Top.scala 31:18]
  wire [15:0] EW_io_Uhht_1_input; // @[Top.scala 31:18]
  wire [15:0] EW_io_output; // @[Top.scala 31:18]
  wire  FC_temp_clock; // @[Top.scala 34:23]
  wire  FC_temp_reset; // @[Top.scala 34:23]
  wire [15:0] FC_temp_io_to_PE_0; // @[Top.scala 34:23]
  wire [15:0] FC_temp_io_to_PE_1; // @[Top.scala 34:23]
  wire [15:0] FC_temp_io_to_PE_2; // @[Top.scala 34:23]
  wire [15:0] FC_temp_io_to_PE_3; // @[Top.scala 34:23]
  wire [15:0] FC_temp_io_to_PE_4; // @[Top.scala 34:23]
  wire [15:0] FC_temp_io_to_PE_5; // @[Top.scala 34:23]
  wire [15:0] FC_temp_io_to_PE_6; // @[Top.scala 34:23]
  wire [15:0] FC_temp_io_to_PE_7; // @[Top.scala 34:23]
  wire [15:0] FC_temp_io_to_PE_8; // @[Top.scala 34:23]
  wire [15:0] FC_temp_io_to_PE_9; // @[Top.scala 34:23]
  wire [15:0] FC_temp_io_to_PE_10; // @[Top.scala 34:23]
  wire [15:0] FC_temp_io_to_PE_11; // @[Top.scala 34:23]
  wire [2:0] FC_temp_io_to_PE_control; // @[Top.scala 34:23]
  wire [15:0] FC_temp_io_rdData; // @[Top.scala 34:23]
  wire  FC_temp_io_wrEna; // @[Top.scala 34:23]
  wire [15:0] FC_temp_io_wrData; // @[Top.scala 34:23]
  wire [5:0] FC_temp_io_wrAddr; // @[Top.scala 34:23]
  wire  Result_clock; // @[Top.scala 35:22]
  wire  Result_reset; // @[Top.scala 35:22]
  wire [15:0] Result_io_rdData; // @[Top.scala 35:22]
  wire  Result_io_wrEna; // @[Top.scala 35:22]
  wire [15:0] Result_io_wrData; // @[Top.scala 35:22]
  wire [3:0] Result_io_wrAddr; // @[Top.scala 35:22]
  wire [15:0] _GEN_12 = FSM_top_io_PE_above_data_ctrl == 2'h2 ? FC_temp_io_to_PE_0 : 16'h0; // @[Top.scala 71:52 Top.scala 72:31 Top.scala 75:36]
  wire [15:0] _GEN_13 = FSM_top_io_PE_above_data_ctrl == 2'h2 ? FC_temp_io_to_PE_1 : 16'h0; // @[Top.scala 71:52 Top.scala 72:31 Top.scala 75:36]
  wire [15:0] _GEN_14 = FSM_top_io_PE_above_data_ctrl == 2'h2 ? FC_temp_io_to_PE_2 : 16'h0; // @[Top.scala 71:52 Top.scala 72:31 Top.scala 75:36]
  wire [15:0] _GEN_15 = FSM_top_io_PE_above_data_ctrl == 2'h2 ? FC_temp_io_to_PE_3 : 16'h0; // @[Top.scala 71:52 Top.scala 72:31 Top.scala 75:36]
  wire [15:0] _GEN_16 = FSM_top_io_PE_above_data_ctrl == 2'h2 ? FC_temp_io_to_PE_4 : 16'h0; // @[Top.scala 71:52 Top.scala 72:31 Top.scala 75:36]
  wire [15:0] _GEN_17 = FSM_top_io_PE_above_data_ctrl == 2'h2 ? FC_temp_io_to_PE_5 : 16'h0; // @[Top.scala 71:52 Top.scala 72:31 Top.scala 75:36]
  wire [15:0] _GEN_18 = FSM_top_io_PE_above_data_ctrl == 2'h2 ? FC_temp_io_to_PE_6 : 16'h0; // @[Top.scala 71:52 Top.scala 72:31 Top.scala 75:36]
  wire [15:0] _GEN_19 = FSM_top_io_PE_above_data_ctrl == 2'h2 ? FC_temp_io_to_PE_7 : 16'h0; // @[Top.scala 71:52 Top.scala 72:31 Top.scala 75:36]
  wire [15:0] _GEN_20 = FSM_top_io_PE_above_data_ctrl == 2'h2 ? FC_temp_io_to_PE_8 : 16'h0; // @[Top.scala 71:52 Top.scala 72:31 Top.scala 75:36]
  wire [15:0] _GEN_21 = FSM_top_io_PE_above_data_ctrl == 2'h2 ? FC_temp_io_to_PE_9 : 16'h0; // @[Top.scala 71:52 Top.scala 72:31 Top.scala 75:36]
  wire [15:0] _GEN_22 = FSM_top_io_PE_above_data_ctrl == 2'h2 ? FC_temp_io_to_PE_10 : 16'h0; // @[Top.scala 71:52 Top.scala 72:31 Top.scala 75:36]
  wire [15:0] _GEN_23 = FSM_top_io_PE_above_data_ctrl == 2'h2 ? FC_temp_io_to_PE_11 : 16'h0; // @[Top.scala 71:52 Top.scala 72:31 Top.scala 75:36]
  wire [15:0] _GEN_24 = FSM_top_io_PE_above_data_ctrl == 2'h1 ? Ht_io_to_PE_0 : _GEN_12; // @[Top.scala 69:52 Top.scala 70:31]
  wire [15:0] _GEN_25 = FSM_top_io_PE_above_data_ctrl == 2'h1 ? Ht_io_to_PE_1 : _GEN_13; // @[Top.scala 69:52 Top.scala 70:31]
  wire [15:0] _GEN_26 = FSM_top_io_PE_above_data_ctrl == 2'h1 ? Ht_io_to_PE_2 : _GEN_14; // @[Top.scala 69:52 Top.scala 70:31]
  wire [15:0] _GEN_27 = FSM_top_io_PE_above_data_ctrl == 2'h1 ? Ht_io_to_PE_3 : _GEN_15; // @[Top.scala 69:52 Top.scala 70:31]
  wire [15:0] _GEN_28 = FSM_top_io_PE_above_data_ctrl == 2'h1 ? Ht_io_to_PE_4 : _GEN_16; // @[Top.scala 69:52 Top.scala 70:31]
  wire [15:0] _GEN_29 = FSM_top_io_PE_above_data_ctrl == 2'h1 ? Ht_io_to_PE_5 : _GEN_17; // @[Top.scala 69:52 Top.scala 70:31]
  wire [15:0] _GEN_30 = FSM_top_io_PE_above_data_ctrl == 2'h1 ? Ht_io_to_PE_6 : _GEN_18; // @[Top.scala 69:52 Top.scala 70:31]
  wire [15:0] _GEN_31 = FSM_top_io_PE_above_data_ctrl == 2'h1 ? Ht_io_to_PE_7 : _GEN_19; // @[Top.scala 69:52 Top.scala 70:31]
  wire [15:0] _GEN_32 = FSM_top_io_PE_above_data_ctrl == 2'h1 ? Ht_io_to_PE_8 : _GEN_20; // @[Top.scala 69:52 Top.scala 70:31]
  wire [15:0] _GEN_33 = FSM_top_io_PE_above_data_ctrl == 2'h1 ? Ht_io_to_PE_9 : _GEN_21; // @[Top.scala 69:52 Top.scala 70:31]
  wire [15:0] _GEN_34 = FSM_top_io_PE_above_data_ctrl == 2'h1 ? Ht_io_to_PE_10 : _GEN_22; // @[Top.scala 69:52 Top.scala 70:31]
  wire [15:0] _GEN_35 = FSM_top_io_PE_above_data_ctrl == 2'h1 ? Ht_io_to_PE_11 : _GEN_23; // @[Top.scala 69:52 Top.scala 70:31]
  Memory L1_Memory_top_0 ( // @[Top.scala 17:42]
    .clock(L1_Memory_top_0_clock),
    .io_rdAddr(L1_Memory_top_0_io_rdAddr),
    .io_rdData(L1_Memory_top_0_io_rdData),
    .io_wrEna(L1_Memory_top_0_io_wrEna),
    .io_wrData(L1_Memory_top_0_io_wrData),
    .io_wrAddr(L1_Memory_top_0_io_wrAddr)
  );
  Memory L1_Memory_top_1 ( // @[Top.scala 17:42]
    .clock(L1_Memory_top_1_clock),
    .io_rdAddr(L1_Memory_top_1_io_rdAddr),
    .io_rdData(L1_Memory_top_1_io_rdData),
    .io_wrEna(L1_Memory_top_1_io_wrEna),
    .io_wrData(L1_Memory_top_1_io_wrData),
    .io_wrAddr(L1_Memory_top_1_io_wrAddr)
  );
  Memory L1_Memory_top_2 ( // @[Top.scala 17:42]
    .clock(L1_Memory_top_2_clock),
    .io_rdAddr(L1_Memory_top_2_io_rdAddr),
    .io_rdData(L1_Memory_top_2_io_rdData),
    .io_wrEna(L1_Memory_top_2_io_wrEna),
    .io_wrData(L1_Memory_top_2_io_wrData),
    .io_wrAddr(L1_Memory_top_2_io_wrAddr)
  );
  Memory L1_Memory_top_3 ( // @[Top.scala 17:42]
    .clock(L1_Memory_top_3_clock),
    .io_rdAddr(L1_Memory_top_3_io_rdAddr),
    .io_rdData(L1_Memory_top_3_io_rdData),
    .io_wrEna(L1_Memory_top_3_io_wrEna),
    .io_wrData(L1_Memory_top_3_io_wrData),
    .io_wrAddr(L1_Memory_top_3_io_wrAddr)
  );
  Memory L1_Memory_top_4 ( // @[Top.scala 17:42]
    .clock(L1_Memory_top_4_clock),
    .io_rdAddr(L1_Memory_top_4_io_rdAddr),
    .io_rdData(L1_Memory_top_4_io_rdData),
    .io_wrEna(L1_Memory_top_4_io_wrEna),
    .io_wrData(L1_Memory_top_4_io_wrData),
    .io_wrAddr(L1_Memory_top_4_io_wrAddr)
  );
  Memory L1_Memory_top_5 ( // @[Top.scala 17:42]
    .clock(L1_Memory_top_5_clock),
    .io_rdAddr(L1_Memory_top_5_io_rdAddr),
    .io_rdData(L1_Memory_top_5_io_rdData),
    .io_wrEna(L1_Memory_top_5_io_wrEna),
    .io_wrData(L1_Memory_top_5_io_wrData),
    .io_wrAddr(L1_Memory_top_5_io_wrAddr)
  );
  Memory L1_Memory_top_6 ( // @[Top.scala 17:42]
    .clock(L1_Memory_top_6_clock),
    .io_rdAddr(L1_Memory_top_6_io_rdAddr),
    .io_rdData(L1_Memory_top_6_io_rdData),
    .io_wrEna(L1_Memory_top_6_io_wrEna),
    .io_wrData(L1_Memory_top_6_io_wrData),
    .io_wrAddr(L1_Memory_top_6_io_wrAddr)
  );
  Memory L1_Memory_top_7 ( // @[Top.scala 17:42]
    .clock(L1_Memory_top_7_clock),
    .io_rdAddr(L1_Memory_top_7_io_rdAddr),
    .io_rdData(L1_Memory_top_7_io_rdData),
    .io_wrEna(L1_Memory_top_7_io_wrEna),
    .io_wrData(L1_Memory_top_7_io_wrData),
    .io_wrAddr(L1_Memory_top_7_io_wrAddr)
  );
  Memory L1_Memory_top_8 ( // @[Top.scala 17:42]
    .clock(L1_Memory_top_8_clock),
    .io_rdAddr(L1_Memory_top_8_io_rdAddr),
    .io_rdData(L1_Memory_top_8_io_rdData),
    .io_wrEna(L1_Memory_top_8_io_wrEna),
    .io_wrData(L1_Memory_top_8_io_wrData),
    .io_wrAddr(L1_Memory_top_8_io_wrAddr)
  );
  Memory L1_Memory_top_9 ( // @[Top.scala 17:42]
    .clock(L1_Memory_top_9_clock),
    .io_rdAddr(L1_Memory_top_9_io_rdAddr),
    .io_rdData(L1_Memory_top_9_io_rdData),
    .io_wrEna(L1_Memory_top_9_io_wrEna),
    .io_wrData(L1_Memory_top_9_io_wrData),
    .io_wrAddr(L1_Memory_top_9_io_wrAddr)
  );
  Memory L1_Memory_top_10 ( // @[Top.scala 17:42]
    .clock(L1_Memory_top_10_clock),
    .io_rdAddr(L1_Memory_top_10_io_rdAddr),
    .io_rdData(L1_Memory_top_10_io_rdData),
    .io_wrEna(L1_Memory_top_10_io_wrEna),
    .io_wrData(L1_Memory_top_10_io_wrData),
    .io_wrAddr(L1_Memory_top_10_io_wrAddr)
  );
  Memory L1_Memory_top_11 ( // @[Top.scala 17:42]
    .clock(L1_Memory_top_11_clock),
    .io_rdAddr(L1_Memory_top_11_io_rdAddr),
    .io_rdData(L1_Memory_top_11_io_rdData),
    .io_wrEna(L1_Memory_top_11_io_wrEna),
    .io_wrData(L1_Memory_top_11_io_wrData),
    .io_wrAddr(L1_Memory_top_11_io_wrAddr)
  );
  PEArray PEArray_top ( // @[Top.scala 18:27]
    .clock(PEArray_top_clock),
    .reset(PEArray_top_reset),
    .io_From_above_0(PEArray_top_io_From_above_0),
    .io_From_above_1(PEArray_top_io_From_above_1),
    .io_From_above_2(PEArray_top_io_From_above_2),
    .io_From_above_3(PEArray_top_io_From_above_3),
    .io_From_above_4(PEArray_top_io_From_above_4),
    .io_From_above_5(PEArray_top_io_From_above_5),
    .io_From_above_6(PEArray_top_io_From_above_6),
    .io_From_above_7(PEArray_top_io_From_above_7),
    .io_From_above_8(PEArray_top_io_From_above_8),
    .io_From_above_9(PEArray_top_io_From_above_9),
    .io_From_above_10(PEArray_top_io_From_above_10),
    .io_From_above_11(PEArray_top_io_From_above_11),
    .io_PE_control_0_mask(PEArray_top_io_PE_control_0_mask),
    .io_PE_control_1_mask(PEArray_top_io_PE_control_1_mask),
    .io_PE_control_2_control(PEArray_top_io_PE_control_2_control),
    .io_PE_control_2_count(PEArray_top_io_PE_control_2_count),
    .io_PE_control_2_L0index(PEArray_top_io_PE_control_2_L0index),
    .io_PE_control_2_mask(PEArray_top_io_PE_control_2_mask),
    .io_PE_control_2_gru_out_width(PEArray_top_io_PE_control_2_gru_out_width),
    .io_rd_data_mux(PEArray_top_io_rd_data_mux),
    .io_To_below_0(PEArray_top_io_To_below_0),
    .io_To_below_1(PEArray_top_io_To_below_1),
    .io_To_below_2(PEArray_top_io_To_below_2),
    .io_To_below_3(PEArray_top_io_To_below_3),
    .io_To_below_4(PEArray_top_io_To_below_4),
    .io_To_below_5(PEArray_top_io_To_below_5),
    .io_To_below_6(PEArray_top_io_To_below_6),
    .io_To_below_7(PEArray_top_io_To_below_7),
    .io_To_below_8(PEArray_top_io_To_below_8),
    .io_To_below_9(PEArray_top_io_To_below_9),
    .io_To_below_10(PEArray_top_io_To_below_10),
    .io_To_below_11(PEArray_top_io_To_below_11),
    .io_To_right_2(PEArray_top_io_To_right_2)
  );
  FSM FSM_top ( // @[Top.scala 19:23]
    .clock(FSM_top_clock),
    .reset(FSM_top_reset),
    .io_Start(FSM_top_io_Start),
    .io_Input_Data(FSM_top_io_Input_Data),
    .io_Input_Valid(FSM_top_io_Input_Valid),
    .io_Input_Ready(FSM_top_io_Input_Ready),
    .io_L1_wr_data(FSM_top_io_L1_wr_data),
    .io_To_L1_control(FSM_top_io_To_L1_control),
    .io_L1_rd_addr_0(FSM_top_io_L1_rd_addr_0),
    .io_L1_rd_addr_1(FSM_top_io_L1_rd_addr_1),
    .io_L1_rd_addr_2(FSM_top_io_L1_rd_addr_2),
    .io_L1_rd_addr_3(FSM_top_io_L1_rd_addr_3),
    .io_L1_rd_addr_4(FSM_top_io_L1_rd_addr_4),
    .io_L1_rd_addr_5(FSM_top_io_L1_rd_addr_5),
    .io_L1_rd_addr_6(FSM_top_io_L1_rd_addr_6),
    .io_L1_rd_addr_7(FSM_top_io_L1_rd_addr_7),
    .io_L1_rd_addr_8(FSM_top_io_L1_rd_addr_8),
    .io_L1_rd_addr_9(FSM_top_io_L1_rd_addr_9),
    .io_L1_rd_addr_10(FSM_top_io_L1_rd_addr_10),
    .io_L1_rd_addr_11(FSM_top_io_L1_rd_addr_11),
    .io_PE_rd_data_mux(FSM_top_io_PE_rd_data_mux),
    .io_L1_wr_addr_0(FSM_top_io_L1_wr_addr_0),
    .io_L1_wr_addr_1(FSM_top_io_L1_wr_addr_1),
    .io_L1_wr_addr_2(FSM_top_io_L1_wr_addr_2),
    .io_L1_wr_addr_3(FSM_top_io_L1_wr_addr_3),
    .io_L1_wr_addr_4(FSM_top_io_L1_wr_addr_4),
    .io_L1_wr_addr_5(FSM_top_io_L1_wr_addr_5),
    .io_L1_wr_addr_6(FSM_top_io_L1_wr_addr_6),
    .io_L1_wr_addr_7(FSM_top_io_L1_wr_addr_7),
    .io_L1_wr_addr_8(FSM_top_io_L1_wr_addr_8),
    .io_L1_wr_addr_9(FSM_top_io_L1_wr_addr_9),
    .io_L1_wr_addr_10(FSM_top_io_L1_wr_addr_10),
    .io_L1_wr_addr_11(FSM_top_io_L1_wr_addr_11),
    .io_L1_wrEna_0(FSM_top_io_L1_wrEna_0),
    .io_L1_wrEna_1(FSM_top_io_L1_wrEna_1),
    .io_L1_wrEna_2(FSM_top_io_L1_wrEna_2),
    .io_L1_wrEna_3(FSM_top_io_L1_wrEna_3),
    .io_L1_wrEna_4(FSM_top_io_L1_wrEna_4),
    .io_L1_wrEna_5(FSM_top_io_L1_wrEna_5),
    .io_L1_wrEna_6(FSM_top_io_L1_wrEna_6),
    .io_L1_wrEna_7(FSM_top_io_L1_wrEna_7),
    .io_L1_wrEna_8(FSM_top_io_L1_wrEna_8),
    .io_L1_wrEna_9(FSM_top_io_L1_wrEna_9),
    .io_L1_wrEna_10(FSM_top_io_L1_wrEna_10),
    .io_L1_wrEna_11(FSM_top_io_L1_wrEna_11),
    .io_PEArray_ctrl_0_mask(FSM_top_io_PEArray_ctrl_0_mask),
    .io_PEArray_ctrl_1_mask(FSM_top_io_PEArray_ctrl_1_mask),
    .io_PEArray_ctrl_2_control(FSM_top_io_PEArray_ctrl_2_control),
    .io_PEArray_ctrl_2_count(FSM_top_io_PEArray_ctrl_2_count),
    .io_PEArray_ctrl_2_L0index(FSM_top_io_PEArray_ctrl_2_L0index),
    .io_PEArray_ctrl_2_mask(FSM_top_io_PEArray_ctrl_2_mask),
    .io_PEArray_ctrl_2_gru_out_width(FSM_top_io_PEArray_ctrl_2_gru_out_width),
    .io_BNArray_ctrl_0(FSM_top_io_BNArray_ctrl_0),
    .io_BNArray_ctrl_1(FSM_top_io_BNArray_ctrl_1),
    .io_BNArray_ctrl_2(FSM_top_io_BNArray_ctrl_2),
    .io_BNArray_ctrl_3(FSM_top_io_BNArray_ctrl_3),
    .io_BNArray_ctrl_4(FSM_top_io_BNArray_ctrl_4),
    .io_BNArray_ctrl_5(FSM_top_io_BNArray_ctrl_5),
    .io_BNArray_ctrl_6(FSM_top_io_BNArray_ctrl_6),
    .io_BNArray_ctrl_7(FSM_top_io_BNArray_ctrl_7),
    .io_BNArray_ctrl_8(FSM_top_io_BNArray_ctrl_8),
    .io_BNArray_ctrl_9(FSM_top_io_BNArray_ctrl_9),
    .io_BNArray_ctrl_10(FSM_top_io_BNArray_ctrl_10),
    .io_BNArray_ctrl_11(FSM_top_io_BNArray_ctrl_11),
    .io_BN_Unit_ctrl(FSM_top_io_BN_Unit_ctrl),
    .io_Relu6Array_ctrl_0(FSM_top_io_Relu6Array_ctrl_0),
    .io_Relu6Array_ctrl_1(FSM_top_io_Relu6Array_ctrl_1),
    .io_Relu6Array_ctrl_2(FSM_top_io_Relu6Array_ctrl_2),
    .io_Relu6Array_ctrl_3(FSM_top_io_Relu6Array_ctrl_3),
    .io_Relu6Array_ctrl_4(FSM_top_io_Relu6Array_ctrl_4),
    .io_Relu6Array_ctrl_5(FSM_top_io_Relu6Array_ctrl_5),
    .io_Relu6Array_ctrl_6(FSM_top_io_Relu6Array_ctrl_6),
    .io_Relu6Array_ctrl_7(FSM_top_io_Relu6Array_ctrl_7),
    .io_Relu6Array_ctrl_8(FSM_top_io_Relu6Array_ctrl_8),
    .io_Relu6Array_ctrl_9(FSM_top_io_Relu6Array_ctrl_9),
    .io_Relu6Array_ctrl_10(FSM_top_io_Relu6Array_ctrl_10),
    .io_Relu6Array_ctrl_11(FSM_top_io_Relu6Array_ctrl_11),
    .io_PE_above_data_ctrl(FSM_top_io_PE_above_data_ctrl),
    .io_Activation_ctrl(FSM_top_io_Activation_ctrl),
    .io_Ht_to_PE_control(FSM_top_io_Ht_to_PE_control),
    .io_Ht_wrEna(FSM_top_io_Ht_wrEna),
    .io_Ht_wrAddr(FSM_top_io_Ht_wrAddr),
    .io_Zt_rdAddr(FSM_top_io_Zt_rdAddr),
    .io_Zt_wrEna(FSM_top_io_Zt_wrEna),
    .io_Zt_wrAddr(FSM_top_io_Zt_wrAddr),
    .io_Rt_rdAddr(FSM_top_io_Rt_rdAddr),
    .io_Rt_wrEna(FSM_top_io_Rt_wrEna),
    .io_Rt_wrAddr(FSM_top_io_Rt_wrAddr),
    .io_WhXt_rdAddr(FSM_top_io_WhXt_rdAddr),
    .io_WhXt_wrEna(FSM_top_io_WhXt_wrEna),
    .io_WhXt_wrAddr(FSM_top_io_WhXt_wrAddr),
    .io_Uhht_1_rdAddr(FSM_top_io_Uhht_1_rdAddr),
    .io_Uhht_1_wrEna(FSM_top_io_Uhht_1_wrEna),
    .io_Uhht_1_wrAddr(FSM_top_io_Uhht_1_wrAddr),
    .io_FC_temp_to_PE_control(FSM_top_io_FC_temp_to_PE_control),
    .io_FC_temp_wrEna(FSM_top_io_FC_temp_wrEna),
    .io_FC_temp_wrAddr(FSM_top_io_FC_temp_wrAddr),
    .io_Result_wrEna(FSM_top_io_Result_wrEna),
    .io_Result_wrAddr(FSM_top_io_Result_wrAddr)
  );
  BN_Unit_Array BN_Array_below ( // @[Top.scala 21:30]
    .clock(BN_Array_below_clock),
    .reset(BN_Array_below_reset),
    .io_from_PE_0(BN_Array_below_io_from_PE_0),
    .io_from_PE_1(BN_Array_below_io_from_PE_1),
    .io_from_PE_2(BN_Array_below_io_from_PE_2),
    .io_from_PE_3(BN_Array_below_io_from_PE_3),
    .io_from_PE_4(BN_Array_below_io_from_PE_4),
    .io_from_PE_5(BN_Array_below_io_from_PE_5),
    .io_from_PE_6(BN_Array_below_io_from_PE_6),
    .io_from_PE_7(BN_Array_below_io_from_PE_7),
    .io_from_PE_8(BN_Array_below_io_from_PE_8),
    .io_from_PE_9(BN_Array_below_io_from_PE_9),
    .io_from_PE_10(BN_Array_below_io_from_PE_10),
    .io_from_PE_11(BN_Array_below_io_from_PE_11),
    .io_control_0(BN_Array_below_io_control_0),
    .io_control_1(BN_Array_below_io_control_1),
    .io_control_2(BN_Array_below_io_control_2),
    .io_control_3(BN_Array_below_io_control_3),
    .io_control_4(BN_Array_below_io_control_4),
    .io_control_5(BN_Array_below_io_control_5),
    .io_control_6(BN_Array_below_io_control_6),
    .io_control_7(BN_Array_below_io_control_7),
    .io_control_8(BN_Array_below_io_control_8),
    .io_control_9(BN_Array_below_io_control_9),
    .io_control_10(BN_Array_below_io_control_10),
    .io_control_11(BN_Array_below_io_control_11),
    .io_to_Relu6_0(BN_Array_below_io_to_Relu6_0),
    .io_to_Relu6_1(BN_Array_below_io_to_Relu6_1),
    .io_to_Relu6_2(BN_Array_below_io_to_Relu6_2),
    .io_to_Relu6_3(BN_Array_below_io_to_Relu6_3),
    .io_to_Relu6_4(BN_Array_below_io_to_Relu6_4),
    .io_to_Relu6_5(BN_Array_below_io_to_Relu6_5),
    .io_to_Relu6_6(BN_Array_below_io_to_Relu6_6),
    .io_to_Relu6_7(BN_Array_below_io_to_Relu6_7),
    .io_to_Relu6_8(BN_Array_below_io_to_Relu6_8),
    .io_to_Relu6_9(BN_Array_below_io_to_Relu6_9),
    .io_to_Relu6_10(BN_Array_below_io_to_Relu6_10),
    .io_to_Relu6_11(BN_Array_below_io_to_Relu6_11)
  );
  Relu6_Unit_Array Relu6_Array ( // @[Top.scala 22:27]
    .io_input_0(Relu6_Array_io_input_0),
    .io_input_1(Relu6_Array_io_input_1),
    .io_input_2(Relu6_Array_io_input_2),
    .io_input_3(Relu6_Array_io_input_3),
    .io_input_4(Relu6_Array_io_input_4),
    .io_input_5(Relu6_Array_io_input_5),
    .io_input_6(Relu6_Array_io_input_6),
    .io_input_7(Relu6_Array_io_input_7),
    .io_input_8(Relu6_Array_io_input_8),
    .io_input_9(Relu6_Array_io_input_9),
    .io_input_10(Relu6_Array_io_input_10),
    .io_input_11(Relu6_Array_io_input_11),
    .io_control_0(Relu6_Array_io_control_0),
    .io_control_1(Relu6_Array_io_control_1),
    .io_control_2(Relu6_Array_io_control_2),
    .io_control_3(Relu6_Array_io_control_3),
    .io_control_4(Relu6_Array_io_control_4),
    .io_control_5(Relu6_Array_io_control_5),
    .io_control_6(Relu6_Array_io_control_6),
    .io_control_7(Relu6_Array_io_control_7),
    .io_control_8(Relu6_Array_io_control_8),
    .io_control_9(Relu6_Array_io_control_9),
    .io_control_10(Relu6_Array_io_control_10),
    .io_control_11(Relu6_Array_io_control_11),
    .io_output_0(Relu6_Array_io_output_0),
    .io_output_1(Relu6_Array_io_output_1),
    .io_output_2(Relu6_Array_io_output_2),
    .io_output_3(Relu6_Array_io_output_3),
    .io_output_4(Relu6_Array_io_output_4),
    .io_output_5(Relu6_Array_io_output_5),
    .io_output_6(Relu6_Array_io_output_6),
    .io_output_7(Relu6_Array_io_output_7),
    .io_output_8(Relu6_Array_io_output_8),
    .io_output_9(Relu6_Array_io_output_9),
    .io_output_10(Relu6_Array_io_output_10),
    .io_output_11(Relu6_Array_io_output_11)
  );
  BN_Unit BNUnit_right ( // @[Top.scala 23:28]
    .clock(BNUnit_right_clock),
    .reset(BNUnit_right_reset),
    .io_input(BNUnit_right_io_input),
    .io_control(BNUnit_right_io_control),
    .io_output(BNUnit_right_io_output)
  );
  activation_Unit Activation ( // @[Top.scala 24:26]
    .clock(Activation_clock),
    .reset(Activation_reset),
    .io_input(Activation_io_input),
    .io_control(Activation_io_control),
    .io_output(Activation_io_output)
  );
  accumulator_registers Zt ( // @[Top.scala 26:18]
    .clock(Zt_clock),
    .reset(Zt_reset),
    .io_rdAddr(Zt_io_rdAddr),
    .io_rdData(Zt_io_rdData),
    .io_wrEna(Zt_io_wrEna),
    .io_wrData(Zt_io_wrData),
    .io_wrAddr(Zt_io_wrAddr)
  );
  accumulator_registers Rt ( // @[Top.scala 27:18]
    .clock(Rt_clock),
    .reset(Rt_reset),
    .io_rdAddr(Rt_io_rdAddr),
    .io_rdData(Rt_io_rdData),
    .io_wrEna(Rt_io_wrEna),
    .io_wrData(Rt_io_wrData),
    .io_wrAddr(Rt_io_wrAddr)
  );
  accumulator_registers WhXt ( // @[Top.scala 28:20]
    .clock(WhXt_clock),
    .reset(WhXt_reset),
    .io_rdAddr(WhXt_io_rdAddr),
    .io_rdData(WhXt_io_rdData),
    .io_wrEna(WhXt_io_wrEna),
    .io_wrData(WhXt_io_wrData),
    .io_wrAddr(WhXt_io_wrAddr)
  );
  accumulator_registers Uhht_1 ( // @[Top.scala 29:22]
    .clock(Uhht_1_clock),
    .reset(Uhht_1_reset),
    .io_rdAddr(Uhht_1_io_rdAddr),
    .io_rdData(Uhht_1_io_rdData),
    .io_wrEna(Uhht_1_io_wrEna),
    .io_wrData(Uhht_1_io_wrData),
    .io_wrAddr(Uhht_1_io_wrAddr)
  );
  ht Ht ( // @[Top.scala 30:18]
    .clock(Ht_clock),
    .reset(Ht_reset),
    .io_to_PE_0(Ht_io_to_PE_0),
    .io_to_PE_1(Ht_io_to_PE_1),
    .io_to_PE_2(Ht_io_to_PE_2),
    .io_to_PE_3(Ht_io_to_PE_3),
    .io_to_PE_4(Ht_io_to_PE_4),
    .io_to_PE_5(Ht_io_to_PE_5),
    .io_to_PE_6(Ht_io_to_PE_6),
    .io_to_PE_7(Ht_io_to_PE_7),
    .io_to_PE_8(Ht_io_to_PE_8),
    .io_to_PE_9(Ht_io_to_PE_9),
    .io_to_PE_10(Ht_io_to_PE_10),
    .io_to_PE_11(Ht_io_to_PE_11),
    .io_to_PE_control(Ht_io_to_PE_control),
    .io_rdData(Ht_io_rdData),
    .io_wrEna(Ht_io_wrEna),
    .io_wrData(Ht_io_wrData),
    .io_wrAddr(Ht_io_wrAddr)
  );
  EW_Unit EW ( // @[Top.scala 31:18]
    .clock(EW_clock),
    .reset(EW_reset),
    .io_ht_1_input(EW_io_ht_1_input),
    .io_Zt_input(EW_io_Zt_input),
    .io_Rt_input(EW_io_Rt_input),
    .io_Whxt_input(EW_io_Whxt_input),
    .io_Uhht_1_input(EW_io_Uhht_1_input),
    .io_output(EW_io_output)
  );
  ht FC_temp ( // @[Top.scala 34:23]
    .clock(FC_temp_clock),
    .reset(FC_temp_reset),
    .io_to_PE_0(FC_temp_io_to_PE_0),
    .io_to_PE_1(FC_temp_io_to_PE_1),
    .io_to_PE_2(FC_temp_io_to_PE_2),
    .io_to_PE_3(FC_temp_io_to_PE_3),
    .io_to_PE_4(FC_temp_io_to_PE_4),
    .io_to_PE_5(FC_temp_io_to_PE_5),
    .io_to_PE_6(FC_temp_io_to_PE_6),
    .io_to_PE_7(FC_temp_io_to_PE_7),
    .io_to_PE_8(FC_temp_io_to_PE_8),
    .io_to_PE_9(FC_temp_io_to_PE_9),
    .io_to_PE_10(FC_temp_io_to_PE_10),
    .io_to_PE_11(FC_temp_io_to_PE_11),
    .io_to_PE_control(FC_temp_io_to_PE_control),
    .io_rdData(FC_temp_io_rdData),
    .io_wrEna(FC_temp_io_wrEna),
    .io_wrData(FC_temp_io_wrData),
    .io_wrAddr(FC_temp_io_wrAddr)
  );
  accumulator_registers_4 Result ( // @[Top.scala 35:22]
    .clock(Result_clock),
    .reset(Result_reset),
    .io_rdData(Result_io_rdData),
    .io_wrEna(Result_io_wrEna),
    .io_wrData(Result_io_wrData),
    .io_wrAddr(Result_io_wrAddr)
  );
  assign io_Input_Ready = 1'h1; // @[Top.scala 151:18]
  assign io_Output_Data = Result_io_rdData; // @[Top.scala 150:18]
  assign L1_Memory_top_0_clock = clock;
  assign L1_Memory_top_0_io_rdAddr = FSM_top_io_L1_rd_addr_0; // @[Top.scala 46:32]
  assign L1_Memory_top_0_io_wrEna = FSM_top_io_L1_wrEna_0; // @[Top.scala 48:32]
  assign L1_Memory_top_0_io_wrData = FSM_top_io_To_L1_control ? FSM_top_io_L1_wr_data : Relu6_Array_io_output_0; // @[Top.scala 51:45 Top.scala 53:34 Top.scala 57:34]
  assign L1_Memory_top_0_io_wrAddr = FSM_top_io_L1_wr_addr_0; // @[Top.scala 47:32]
  assign L1_Memory_top_1_clock = clock;
  assign L1_Memory_top_1_io_rdAddr = FSM_top_io_L1_rd_addr_1; // @[Top.scala 46:32]
  assign L1_Memory_top_1_io_wrEna = FSM_top_io_L1_wrEna_1; // @[Top.scala 48:32]
  assign L1_Memory_top_1_io_wrData = FSM_top_io_To_L1_control ? FSM_top_io_L1_wr_data : Relu6_Array_io_output_1; // @[Top.scala 51:45 Top.scala 53:34 Top.scala 57:34]
  assign L1_Memory_top_1_io_wrAddr = FSM_top_io_L1_wr_addr_1; // @[Top.scala 47:32]
  assign L1_Memory_top_2_clock = clock;
  assign L1_Memory_top_2_io_rdAddr = FSM_top_io_L1_rd_addr_2; // @[Top.scala 46:32]
  assign L1_Memory_top_2_io_wrEna = FSM_top_io_L1_wrEna_2; // @[Top.scala 48:32]
  assign L1_Memory_top_2_io_wrData = FSM_top_io_To_L1_control ? FSM_top_io_L1_wr_data : Relu6_Array_io_output_2; // @[Top.scala 51:45 Top.scala 53:34 Top.scala 57:34]
  assign L1_Memory_top_2_io_wrAddr = FSM_top_io_L1_wr_addr_2; // @[Top.scala 47:32]
  assign L1_Memory_top_3_clock = clock;
  assign L1_Memory_top_3_io_rdAddr = FSM_top_io_L1_rd_addr_3; // @[Top.scala 46:32]
  assign L1_Memory_top_3_io_wrEna = FSM_top_io_L1_wrEna_3; // @[Top.scala 48:32]
  assign L1_Memory_top_3_io_wrData = FSM_top_io_To_L1_control ? FSM_top_io_L1_wr_data : Relu6_Array_io_output_3; // @[Top.scala 51:45 Top.scala 53:34 Top.scala 57:34]
  assign L1_Memory_top_3_io_wrAddr = FSM_top_io_L1_wr_addr_3; // @[Top.scala 47:32]
  assign L1_Memory_top_4_clock = clock;
  assign L1_Memory_top_4_io_rdAddr = FSM_top_io_L1_rd_addr_4; // @[Top.scala 46:32]
  assign L1_Memory_top_4_io_wrEna = FSM_top_io_L1_wrEna_4; // @[Top.scala 48:32]
  assign L1_Memory_top_4_io_wrData = FSM_top_io_To_L1_control ? FSM_top_io_L1_wr_data : Relu6_Array_io_output_4; // @[Top.scala 51:45 Top.scala 53:34 Top.scala 57:34]
  assign L1_Memory_top_4_io_wrAddr = FSM_top_io_L1_wr_addr_4; // @[Top.scala 47:32]
  assign L1_Memory_top_5_clock = clock;
  assign L1_Memory_top_5_io_rdAddr = FSM_top_io_L1_rd_addr_5; // @[Top.scala 46:32]
  assign L1_Memory_top_5_io_wrEna = FSM_top_io_L1_wrEna_5; // @[Top.scala 48:32]
  assign L1_Memory_top_5_io_wrData = FSM_top_io_To_L1_control ? FSM_top_io_L1_wr_data : Relu6_Array_io_output_5; // @[Top.scala 51:45 Top.scala 53:34 Top.scala 57:34]
  assign L1_Memory_top_5_io_wrAddr = FSM_top_io_L1_wr_addr_5; // @[Top.scala 47:32]
  assign L1_Memory_top_6_clock = clock;
  assign L1_Memory_top_6_io_rdAddr = FSM_top_io_L1_rd_addr_6; // @[Top.scala 46:32]
  assign L1_Memory_top_6_io_wrEna = FSM_top_io_L1_wrEna_6; // @[Top.scala 48:32]
  assign L1_Memory_top_6_io_wrData = FSM_top_io_To_L1_control ? FSM_top_io_L1_wr_data : Relu6_Array_io_output_6; // @[Top.scala 51:45 Top.scala 53:34 Top.scala 57:34]
  assign L1_Memory_top_6_io_wrAddr = FSM_top_io_L1_wr_addr_6; // @[Top.scala 47:32]
  assign L1_Memory_top_7_clock = clock;
  assign L1_Memory_top_7_io_rdAddr = FSM_top_io_L1_rd_addr_7; // @[Top.scala 46:32]
  assign L1_Memory_top_7_io_wrEna = FSM_top_io_L1_wrEna_7; // @[Top.scala 48:32]
  assign L1_Memory_top_7_io_wrData = FSM_top_io_To_L1_control ? FSM_top_io_L1_wr_data : Relu6_Array_io_output_7; // @[Top.scala 51:45 Top.scala 53:34 Top.scala 57:34]
  assign L1_Memory_top_7_io_wrAddr = FSM_top_io_L1_wr_addr_7; // @[Top.scala 47:32]
  assign L1_Memory_top_8_clock = clock;
  assign L1_Memory_top_8_io_rdAddr = FSM_top_io_L1_rd_addr_8; // @[Top.scala 46:32]
  assign L1_Memory_top_8_io_wrEna = FSM_top_io_L1_wrEna_8; // @[Top.scala 48:32]
  assign L1_Memory_top_8_io_wrData = FSM_top_io_To_L1_control ? FSM_top_io_L1_wr_data : Relu6_Array_io_output_8; // @[Top.scala 51:45 Top.scala 53:34 Top.scala 57:34]
  assign L1_Memory_top_8_io_wrAddr = FSM_top_io_L1_wr_addr_8; // @[Top.scala 47:32]
  assign L1_Memory_top_9_clock = clock;
  assign L1_Memory_top_9_io_rdAddr = FSM_top_io_L1_rd_addr_9; // @[Top.scala 46:32]
  assign L1_Memory_top_9_io_wrEna = FSM_top_io_L1_wrEna_9; // @[Top.scala 48:32]
  assign L1_Memory_top_9_io_wrData = FSM_top_io_To_L1_control ? FSM_top_io_L1_wr_data : Relu6_Array_io_output_9; // @[Top.scala 51:45 Top.scala 53:34 Top.scala 57:34]
  assign L1_Memory_top_9_io_wrAddr = FSM_top_io_L1_wr_addr_9; // @[Top.scala 47:32]
  assign L1_Memory_top_10_clock = clock;
  assign L1_Memory_top_10_io_rdAddr = FSM_top_io_L1_rd_addr_10; // @[Top.scala 46:32]
  assign L1_Memory_top_10_io_wrEna = FSM_top_io_L1_wrEna_10; // @[Top.scala 48:32]
  assign L1_Memory_top_10_io_wrData = FSM_top_io_To_L1_control ? FSM_top_io_L1_wr_data : Relu6_Array_io_output_10; // @[Top.scala 51:45 Top.scala 53:34 Top.scala 57:34]
  assign L1_Memory_top_10_io_wrAddr = FSM_top_io_L1_wr_addr_10; // @[Top.scala 47:32]
  assign L1_Memory_top_11_clock = clock;
  assign L1_Memory_top_11_io_rdAddr = FSM_top_io_L1_rd_addr_11; // @[Top.scala 46:32]
  assign L1_Memory_top_11_io_wrEna = FSM_top_io_L1_wrEna_11; // @[Top.scala 48:32]
  assign L1_Memory_top_11_io_wrData = FSM_top_io_To_L1_control ? FSM_top_io_L1_wr_data : Relu6_Array_io_output_11; // @[Top.scala 51:45 Top.scala 53:34 Top.scala 57:34]
  assign L1_Memory_top_11_io_wrAddr = FSM_top_io_L1_wr_addr_11; // @[Top.scala 47:32]
  assign PEArray_top_clock = clock;
  assign PEArray_top_reset = reset;
  assign PEArray_top_io_From_above_0 = FSM_top_io_PE_above_data_ctrl == 2'h0 ? L1_Memory_top_0_io_rdData : _GEN_24; // @[Top.scala 65:46 Top.scala 67:36]
  assign PEArray_top_io_From_above_1 = FSM_top_io_PE_above_data_ctrl == 2'h0 ? L1_Memory_top_1_io_rdData : _GEN_25; // @[Top.scala 65:46 Top.scala 67:36]
  assign PEArray_top_io_From_above_2 = FSM_top_io_PE_above_data_ctrl == 2'h0 ? L1_Memory_top_2_io_rdData : _GEN_26; // @[Top.scala 65:46 Top.scala 67:36]
  assign PEArray_top_io_From_above_3 = FSM_top_io_PE_above_data_ctrl == 2'h0 ? L1_Memory_top_3_io_rdData : _GEN_27; // @[Top.scala 65:46 Top.scala 67:36]
  assign PEArray_top_io_From_above_4 = FSM_top_io_PE_above_data_ctrl == 2'h0 ? L1_Memory_top_4_io_rdData : _GEN_28; // @[Top.scala 65:46 Top.scala 67:36]
  assign PEArray_top_io_From_above_5 = FSM_top_io_PE_above_data_ctrl == 2'h0 ? L1_Memory_top_5_io_rdData : _GEN_29; // @[Top.scala 65:46 Top.scala 67:36]
  assign PEArray_top_io_From_above_6 = FSM_top_io_PE_above_data_ctrl == 2'h0 ? L1_Memory_top_6_io_rdData : _GEN_30; // @[Top.scala 65:46 Top.scala 67:36]
  assign PEArray_top_io_From_above_7 = FSM_top_io_PE_above_data_ctrl == 2'h0 ? L1_Memory_top_7_io_rdData : _GEN_31; // @[Top.scala 65:46 Top.scala 67:36]
  assign PEArray_top_io_From_above_8 = FSM_top_io_PE_above_data_ctrl == 2'h0 ? L1_Memory_top_8_io_rdData : _GEN_32; // @[Top.scala 65:46 Top.scala 67:36]
  assign PEArray_top_io_From_above_9 = FSM_top_io_PE_above_data_ctrl == 2'h0 ? L1_Memory_top_9_io_rdData : _GEN_33; // @[Top.scala 65:46 Top.scala 67:36]
  assign PEArray_top_io_From_above_10 = FSM_top_io_PE_above_data_ctrl == 2'h0 ? L1_Memory_top_10_io_rdData : _GEN_34; // @[Top.scala 65:46 Top.scala 67:36]
  assign PEArray_top_io_From_above_11 = FSM_top_io_PE_above_data_ctrl == 2'h0 ? L1_Memory_top_11_io_rdData : _GEN_35; // @[Top.scala 65:46 Top.scala 67:36]
  assign PEArray_top_io_PE_control_0_mask = FSM_top_io_PEArray_ctrl_0_mask; // @[Top.scala 62:31]
  assign PEArray_top_io_PE_control_1_mask = FSM_top_io_PEArray_ctrl_1_mask; // @[Top.scala 62:31]
  assign PEArray_top_io_PE_control_2_control = FSM_top_io_PEArray_ctrl_2_control; // @[Top.scala 62:31]
  assign PEArray_top_io_PE_control_2_count = FSM_top_io_PEArray_ctrl_2_count; // @[Top.scala 62:31]
  assign PEArray_top_io_PE_control_2_L0index = FSM_top_io_PEArray_ctrl_2_L0index; // @[Top.scala 62:31]
  assign PEArray_top_io_PE_control_2_mask = FSM_top_io_PEArray_ctrl_2_mask; // @[Top.scala 62:31]
  assign PEArray_top_io_PE_control_2_gru_out_width = FSM_top_io_PEArray_ctrl_2_gru_out_width; // @[Top.scala 62:31]
  assign PEArray_top_io_rd_data_mux = FSM_top_io_PE_rd_data_mux; // @[Top.scala 63:31]
  assign FSM_top_clock = clock;
  assign FSM_top_reset = reset;
  assign FSM_top_io_Start = io_Start; // @[Top.scala 39:21]
  assign FSM_top_io_Input_Data = io_Input_Data; // @[Top.scala 40:27]
  assign FSM_top_io_Input_Valid = io_Input_Valid; // @[Top.scala 41:27]
  assign BN_Array_below_clock = clock;
  assign BN_Array_below_reset = reset;
  assign BN_Array_below_io_from_PE_0 = PEArray_top_io_To_below_0; // @[Top.scala 82:29]
  assign BN_Array_below_io_from_PE_1 = PEArray_top_io_To_below_1; // @[Top.scala 82:29]
  assign BN_Array_below_io_from_PE_2 = PEArray_top_io_To_below_2; // @[Top.scala 82:29]
  assign BN_Array_below_io_from_PE_3 = PEArray_top_io_To_below_3; // @[Top.scala 82:29]
  assign BN_Array_below_io_from_PE_4 = PEArray_top_io_To_below_4; // @[Top.scala 82:29]
  assign BN_Array_below_io_from_PE_5 = PEArray_top_io_To_below_5; // @[Top.scala 82:29]
  assign BN_Array_below_io_from_PE_6 = PEArray_top_io_To_below_6; // @[Top.scala 82:29]
  assign BN_Array_below_io_from_PE_7 = PEArray_top_io_To_below_7; // @[Top.scala 82:29]
  assign BN_Array_below_io_from_PE_8 = PEArray_top_io_To_below_8; // @[Top.scala 82:29]
  assign BN_Array_below_io_from_PE_9 = PEArray_top_io_To_below_9; // @[Top.scala 82:29]
  assign BN_Array_below_io_from_PE_10 = PEArray_top_io_To_below_10; // @[Top.scala 82:29]
  assign BN_Array_below_io_from_PE_11 = PEArray_top_io_To_below_11; // @[Top.scala 82:29]
  assign BN_Array_below_io_control_0 = FSM_top_io_BNArray_ctrl_0; // @[Top.scala 81:29]
  assign BN_Array_below_io_control_1 = FSM_top_io_BNArray_ctrl_1; // @[Top.scala 81:29]
  assign BN_Array_below_io_control_2 = FSM_top_io_BNArray_ctrl_2; // @[Top.scala 81:29]
  assign BN_Array_below_io_control_3 = FSM_top_io_BNArray_ctrl_3; // @[Top.scala 81:29]
  assign BN_Array_below_io_control_4 = FSM_top_io_BNArray_ctrl_4; // @[Top.scala 81:29]
  assign BN_Array_below_io_control_5 = FSM_top_io_BNArray_ctrl_5; // @[Top.scala 81:29]
  assign BN_Array_below_io_control_6 = FSM_top_io_BNArray_ctrl_6; // @[Top.scala 81:29]
  assign BN_Array_below_io_control_7 = FSM_top_io_BNArray_ctrl_7; // @[Top.scala 81:29]
  assign BN_Array_below_io_control_8 = FSM_top_io_BNArray_ctrl_8; // @[Top.scala 81:29]
  assign BN_Array_below_io_control_9 = FSM_top_io_BNArray_ctrl_9; // @[Top.scala 81:29]
  assign BN_Array_below_io_control_10 = FSM_top_io_BNArray_ctrl_10; // @[Top.scala 81:29]
  assign BN_Array_below_io_control_11 = FSM_top_io_BNArray_ctrl_11; // @[Top.scala 81:29]
  assign Relu6_Array_io_input_0 = BN_Array_below_io_to_Relu6_0; // @[Top.scala 96:24]
  assign Relu6_Array_io_input_1 = BN_Array_below_io_to_Relu6_1; // @[Top.scala 96:24]
  assign Relu6_Array_io_input_2 = BN_Array_below_io_to_Relu6_2; // @[Top.scala 96:24]
  assign Relu6_Array_io_input_3 = BN_Array_below_io_to_Relu6_3; // @[Top.scala 96:24]
  assign Relu6_Array_io_input_4 = BN_Array_below_io_to_Relu6_4; // @[Top.scala 96:24]
  assign Relu6_Array_io_input_5 = BN_Array_below_io_to_Relu6_5; // @[Top.scala 96:24]
  assign Relu6_Array_io_input_6 = BN_Array_below_io_to_Relu6_6; // @[Top.scala 96:24]
  assign Relu6_Array_io_input_7 = BN_Array_below_io_to_Relu6_7; // @[Top.scala 96:24]
  assign Relu6_Array_io_input_8 = BN_Array_below_io_to_Relu6_8; // @[Top.scala 96:24]
  assign Relu6_Array_io_input_9 = BN_Array_below_io_to_Relu6_9; // @[Top.scala 96:24]
  assign Relu6_Array_io_input_10 = BN_Array_below_io_to_Relu6_10; // @[Top.scala 96:24]
  assign Relu6_Array_io_input_11 = BN_Array_below_io_to_Relu6_11; // @[Top.scala 96:24]
  assign Relu6_Array_io_control_0 = FSM_top_io_Relu6Array_ctrl_0; // @[Top.scala 95:26]
  assign Relu6_Array_io_control_1 = FSM_top_io_Relu6Array_ctrl_1; // @[Top.scala 95:26]
  assign Relu6_Array_io_control_2 = FSM_top_io_Relu6Array_ctrl_2; // @[Top.scala 95:26]
  assign Relu6_Array_io_control_3 = FSM_top_io_Relu6Array_ctrl_3; // @[Top.scala 95:26]
  assign Relu6_Array_io_control_4 = FSM_top_io_Relu6Array_ctrl_4; // @[Top.scala 95:26]
  assign Relu6_Array_io_control_5 = FSM_top_io_Relu6Array_ctrl_5; // @[Top.scala 95:26]
  assign Relu6_Array_io_control_6 = FSM_top_io_Relu6Array_ctrl_6; // @[Top.scala 95:26]
  assign Relu6_Array_io_control_7 = FSM_top_io_Relu6Array_ctrl_7; // @[Top.scala 95:26]
  assign Relu6_Array_io_control_8 = FSM_top_io_Relu6Array_ctrl_8; // @[Top.scala 95:26]
  assign Relu6_Array_io_control_9 = FSM_top_io_Relu6Array_ctrl_9; // @[Top.scala 95:26]
  assign Relu6_Array_io_control_10 = FSM_top_io_Relu6Array_ctrl_10; // @[Top.scala 95:26]
  assign Relu6_Array_io_control_11 = FSM_top_io_Relu6Array_ctrl_11; // @[Top.scala 95:26]
  assign BNUnit_right_clock = clock;
  assign BNUnit_right_reset = reset;
  assign BNUnit_right_io_input = PEArray_top_io_To_right_2; // @[Top.scala 89:29]
  assign BNUnit_right_io_control = FSM_top_io_BN_Unit_ctrl; // @[Top.scala 88:29]
  assign Activation_clock = clock;
  assign Activation_reset = reset;
  assign Activation_io_input = BNUnit_right_io_output; // @[Top.scala 99:25]
  assign Activation_io_control = FSM_top_io_Activation_ctrl; // @[Top.scala 100:25]
  assign Zt_clock = clock;
  assign Zt_reset = reset;
  assign Zt_io_rdAddr = FSM_top_io_Zt_rdAddr; // @[Top.scala 112:17]
  assign Zt_io_wrEna = FSM_top_io_Zt_wrEna; // @[Top.scala 110:17]
  assign Zt_io_wrData = Activation_io_output; // @[Top.scala 109:17]
  assign Zt_io_wrAddr = FSM_top_io_Zt_wrAddr; // @[Top.scala 111:17]
  assign Rt_clock = clock;
  assign Rt_reset = reset;
  assign Rt_io_rdAddr = FSM_top_io_Rt_rdAddr; // @[Top.scala 117:17]
  assign Rt_io_wrEna = FSM_top_io_Rt_wrEna; // @[Top.scala 115:17]
  assign Rt_io_wrData = Activation_io_output; // @[Top.scala 114:17]
  assign Rt_io_wrAddr = FSM_top_io_Rt_wrAddr; // @[Top.scala 116:17]
  assign WhXt_clock = clock;
  assign WhXt_reset = reset;
  assign WhXt_io_rdAddr = FSM_top_io_WhXt_rdAddr; // @[Top.scala 122:19]
  assign WhXt_io_wrEna = FSM_top_io_WhXt_wrEna; // @[Top.scala 120:19]
  assign WhXt_io_wrData = Activation_io_output; // @[Top.scala 119:19]
  assign WhXt_io_wrAddr = FSM_top_io_WhXt_wrAddr; // @[Top.scala 121:19]
  assign Uhht_1_clock = clock;
  assign Uhht_1_reset = reset;
  assign Uhht_1_io_rdAddr = FSM_top_io_Uhht_1_rdAddr; // @[Top.scala 127:21]
  assign Uhht_1_io_wrEna = FSM_top_io_Uhht_1_wrEna; // @[Top.scala 125:21]
  assign Uhht_1_io_wrData = Activation_io_output; // @[Top.scala 124:21]
  assign Uhht_1_io_wrAddr = FSM_top_io_Uhht_1_wrAddr; // @[Top.scala 126:21]
  assign Ht_clock = clock;
  assign Ht_reset = reset;
  assign Ht_io_to_PE_control = FSM_top_io_Ht_to_PE_control; // @[Top.scala 107:23]
  assign Ht_io_wrEna = FSM_top_io_Ht_wrEna; // @[Top.scala 104:23]
  assign Ht_io_wrData = EW_io_output; // @[Top.scala 103:23]
  assign Ht_io_wrAddr = FSM_top_io_Ht_wrAddr; // @[Top.scala 105:23]
  assign EW_clock = clock;
  assign EW_reset = reset;
  assign EW_io_ht_1_input = Ht_io_rdData; // @[Top.scala 130:23]
  assign EW_io_Zt_input = Zt_io_rdData; // @[Top.scala 131:23]
  assign EW_io_Rt_input = Rt_io_rdData; // @[Top.scala 132:23]
  assign EW_io_Whxt_input = WhXt_io_rdData; // @[Top.scala 133:23]
  assign EW_io_Uhht_1_input = Uhht_1_io_rdData; // @[Top.scala 134:23]
  assign FC_temp_clock = clock;
  assign FC_temp_reset = reset;
  assign FC_temp_io_to_PE_control = FSM_top_io_FC_temp_to_PE_control; // @[Top.scala 141:28]
  assign FC_temp_io_wrEna = FSM_top_io_FC_temp_wrEna; // @[Top.scala 138:28]
  assign FC_temp_io_wrData = Activation_io_output; // @[Top.scala 137:28]
  assign FC_temp_io_wrAddr = FSM_top_io_FC_temp_wrAddr; // @[Top.scala 139:28]
  assign Result_clock = clock;
  assign Result_reset = reset;
  assign Result_io_wrEna = FSM_top_io_Result_wrEna; // @[Top.scala 145:21]
  assign Result_io_wrData = Activation_io_output; // @[Top.scala 144:21]
  assign Result_io_wrAddr = FSM_top_io_Result_wrAddr; // @[Top.scala 146:21]
endmodule
